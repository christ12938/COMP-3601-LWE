----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/16/2021 04:58:20 PM
-- Design Name: 
-- Module Name: log_deltas - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE WORK.DATA_TYPES.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity exp_deltas is
    Port (frac : in unsigned(10 downto 0);
          delta : out unsigned(k_trunc-1 downto 0));
end exp_deltas;

architecture Behavioral of exp_deltas is
begin

process (frac)
begin
    case frac is
        when "00000000000" => delta <= "000000000000010";
        when "00000000001" => delta <= "000000000000111";
        when "00000000010" => delta <= "000000000001100";
        when "00000000011" => delta <= "000000000010001";
        when "00000000100" => delta <= "000000000010101";
        when "00000000101" => delta <= "000000000011010";
        when "00000000110" => delta <= "000000000011111";
        when "00000000111" => delta <= "000000000100100";
        when "00000001000" => delta <= "000000000101001";
        when "00000001001" => delta <= "000000000101110";
        when "00000001010" => delta <= "000000000110011";
        when "00000001011" => delta <= "000000000111000";
        when "00000001100" => delta <= "000000000111100";
        when "00000001101" => delta <= "000000001000001";
        when "00000001110" => delta <= "000000001000110";
        when "00000001111" => delta <= "000000001001011";
        when "00000010000" => delta <= "000000001010000";
        when "00000010001" => delta <= "000000001010101";
        when "00000010010" => delta <= "000000001011010";
        when "00000010011" => delta <= "000000001011110";
        when "00000010100" => delta <= "000000001100011";
        when "00000010101" => delta <= "000000001101000";
        when "00000010110" => delta <= "000000001101101";
        when "00000010111" => delta <= "000000001110010";
        when "00000011000" => delta <= "000000001110111";
        when "00000011001" => delta <= "000000001111011";
        when "00000011010" => delta <= "000000010000000";
        when "00000011011" => delta <= "000000010000101";
        when "00000011100" => delta <= "000000010001010";
        when "00000011101" => delta <= "000000010001111";
        when "00000011110" => delta <= "000000010010011";
        when "00000011111" => delta <= "000000010011000";
        when "00000100000" => delta <= "000000010011101";
        when "00000100001" => delta <= "000000010100010";
        when "00000100010" => delta <= "000000010100110";
        when "00000100011" => delta <= "000000010101011";
        when "00000100100" => delta <= "000000010110000";
        when "00000100101" => delta <= "000000010110101";
        when "00000100110" => delta <= "000000010111010";
        when "00000100111" => delta <= "000000010111110";
        when "00000101000" => delta <= "000000011000011";
        when "00000101001" => delta <= "000000011001000";
        when "00000101010" => delta <= "000000011001101";
        when "00000101011" => delta <= "000000011010001";
        when "00000101100" => delta <= "000000011010110";
        when "00000101101" => delta <= "000000011011011";
        when "00000101110" => delta <= "000000011100000";
        when "00000101111" => delta <= "000000011100100";
        when "00000110000" => delta <= "000000011101001";
        when "00000110001" => delta <= "000000011101110";
        when "00000110010" => delta <= "000000011110010";
        when "00000110011" => delta <= "000000011110111";
        when "00000110100" => delta <= "000000011111100";
        when "00000110101" => delta <= "000000100000001";
        when "00000110110" => delta <= "000000100000101";
        when "00000110111" => delta <= "000000100001010";
        when "00000111000" => delta <= "000000100001111";
        when "00000111001" => delta <= "000000100010011";
        when "00000111010" => delta <= "000000100011000";
        when "00000111011" => delta <= "000000100011101";
        when "00000111100" => delta <= "000000100100001";
        when "00000111101" => delta <= "000000100100110";
        when "00000111110" => delta <= "000000100101011";
        when "00000111111" => delta <= "000000100101111";
        when "00001000000" => delta <= "000000100110100";
        when "00001000001" => delta <= "000000100111001";
        when "00001000010" => delta <= "000000100111101";
        when "00001000011" => delta <= "000000101000010";
        when "00001000100" => delta <= "000000101000111";
        when "00001000101" => delta <= "000000101001011";
        when "00001000110" => delta <= "000000101010000";
        when "00001000111" => delta <= "000000101010101";
        when "00001001000" => delta <= "000000101011001";
        when "00001001001" => delta <= "000000101011110";
        when "00001001010" => delta <= "000000101100011";
        when "00001001011" => delta <= "000000101100111";
        when "00001001100" => delta <= "000000101101100";
        when "00001001101" => delta <= "000000101110000";
        when "00001001110" => delta <= "000000101110101";
        when "00001001111" => delta <= "000000101111010";
        when "00001010000" => delta <= "000000101111110";
        when "00001010001" => delta <= "000000110000011";
        when "00001010010" => delta <= "000000110001000";
        when "00001010011" => delta <= "000000110001100";
        when "00001010100" => delta <= "000000110010001";
        when "00001010101" => delta <= "000000110010101";
        when "00001010110" => delta <= "000000110011010";
        when "00001010111" => delta <= "000000110011110";
        when "00001011000" => delta <= "000000110100011";
        when "00001011001" => delta <= "000000110101000";
        when "00001011010" => delta <= "000000110101100";
        when "00001011011" => delta <= "000000110110001";
        when "00001011100" => delta <= "000000110110101";
        when "00001011101" => delta <= "000000110111010";
        when "00001011110" => delta <= "000000110111110";
        when "00001011111" => delta <= "000000111000011";
        when "00001100000" => delta <= "000000111000111";
        when "00001100001" => delta <= "000000111001100";
        when "00001100010" => delta <= "000000111010001";
        when "00001100011" => delta <= "000000111010101";
        when "00001100100" => delta <= "000000111011010";
        when "00001100101" => delta <= "000000111011110";
        when "00001100110" => delta <= "000000111100011";
        when "00001100111" => delta <= "000000111100111";
        when "00001101000" => delta <= "000000111101100";
        when "00001101001" => delta <= "000000111110000";
        when "00001101010" => delta <= "000000111110101";
        when "00001101011" => delta <= "000000111111001";
        when "00001101100" => delta <= "000000111111110";
        when "00001101101" => delta <= "000001000000010";
        when "00001101110" => delta <= "000001000000111";
        when "00001101111" => delta <= "000001000001011";
        when "00001110000" => delta <= "000001000010000";
        when "00001110001" => delta <= "000001000010100";
        when "00001110010" => delta <= "000001000011001";
        when "00001110011" => delta <= "000001000011101";
        when "00001110100" => delta <= "000001000100010";
        when "00001110101" => delta <= "000001000100110";
        when "00001110110" => delta <= "000001000101010";
        when "00001110111" => delta <= "000001000101111";
        when "00001111000" => delta <= "000001000110011";
        when "00001111001" => delta <= "000001000111000";
        when "00001111010" => delta <= "000001000111100";
        when "00001111011" => delta <= "000001001000001";
        when "00001111100" => delta <= "000001001000101";
        when "00001111101" => delta <= "000001001001010";
        when "00001111110" => delta <= "000001001001110";
        when "00001111111" => delta <= "000001001010010";
        when "00010000000" => delta <= "000001001010111";
        when "00010000001" => delta <= "000001001011011";
        when "00010000010" => delta <= "000001001100000";
        when "00010000011" => delta <= "000001001100100";
        when "00010000100" => delta <= "000001001101000";
        when "00010000101" => delta <= "000001001101101";
        when "00010000110" => delta <= "000001001110001";
        when "00010000111" => delta <= "000001001110110";
        when "00010001000" => delta <= "000001001111010";
        when "00010001001" => delta <= "000001001111110";
        when "00010001010" => delta <= "000001010000011";
        when "00010001011" => delta <= "000001010000111";
        when "00010001100" => delta <= "000001010001100";
        when "00010001101" => delta <= "000001010010000";
        when "00010001110" => delta <= "000001010010100";
        when "00010001111" => delta <= "000001010011001";
        when "00010010000" => delta <= "000001010011101";
        when "00010010001" => delta <= "000001010100001";
        when "00010010010" => delta <= "000001010100110";
        when "00010010011" => delta <= "000001010101010";
        when "00010010100" => delta <= "000001010101110";
        when "00010010101" => delta <= "000001010110011";
        when "00010010110" => delta <= "000001010110111";
        when "00010010111" => delta <= "000001010111011";
        when "00010011000" => delta <= "000001011000000";
        when "00010011001" => delta <= "000001011000100";
        when "00010011010" => delta <= "000001011001000";
        when "00010011011" => delta <= "000001011001101";
        when "00010011100" => delta <= "000001011010001";
        when "00010011101" => delta <= "000001011010101";
        when "00010011110" => delta <= "000001011011010";
        when "00010011111" => delta <= "000001011011110";
        when "00010100000" => delta <= "000001011100010";
        when "00010100001" => delta <= "000001011100110";
        when "00010100010" => delta <= "000001011101011";
        when "00010100011" => delta <= "000001011101111";
        when "00010100100" => delta <= "000001011110011";
        when "00010100101" => delta <= "000001011111000";
        when "00010100110" => delta <= "000001011111100";
        when "00010100111" => delta <= "000001100000000";
        when "00010101000" => delta <= "000001100000100";
        when "00010101001" => delta <= "000001100001001";
        when "00010101010" => delta <= "000001100001101";
        when "00010101011" => delta <= "000001100010001";
        when "00010101100" => delta <= "000001100010101";
        when "00010101101" => delta <= "000001100011010";
        when "00010101110" => delta <= "000001100011110";
        when "00010101111" => delta <= "000001100100010";
        when "00010110000" => delta <= "000001100100110";
        when "00010110001" => delta <= "000001100101010";
        when "00010110010" => delta <= "000001100101111";
        when "00010110011" => delta <= "000001100110011";
        when "00010110100" => delta <= "000001100110111";
        when "00010110101" => delta <= "000001100111011";
        when "00010110110" => delta <= "000001101000000";
        when "00010110111" => delta <= "000001101000100";
        when "00010111000" => delta <= "000001101001000";
        when "00010111001" => delta <= "000001101001100";
        when "00010111010" => delta <= "000001101010000";
        when "00010111011" => delta <= "000001101010101";
        when "00010111100" => delta <= "000001101011001";
        when "00010111101" => delta <= "000001101011101";
        when "00010111110" => delta <= "000001101100001";
        when "00010111111" => delta <= "000001101100101";
        when "00011000000" => delta <= "000001101101001";
        when "00011000001" => delta <= "000001101101110";
        when "00011000010" => delta <= "000001101110010";
        when "00011000011" => delta <= "000001101110110";
        when "00011000100" => delta <= "000001101111010";
        when "00011000101" => delta <= "000001101111110";
        when "00011000110" => delta <= "000001110000010";
        when "00011000111" => delta <= "000001110000110";
        when "00011001000" => delta <= "000001110001011";
        when "00011001001" => delta <= "000001110001111";
        when "00011001010" => delta <= "000001110010011";
        when "00011001011" => delta <= "000001110010111";
        when "00011001100" => delta <= "000001110011011";
        when "00011001101" => delta <= "000001110011111";
        when "00011001110" => delta <= "000001110100011";
        when "00011001111" => delta <= "000001110100111";
        when "00011010000" => delta <= "000001110101011";
        when "00011010001" => delta <= "000001110110000";
        when "00011010010" => delta <= "000001110110100";
        when "00011010011" => delta <= "000001110111000";
        when "00011010100" => delta <= "000001110111100";
        when "00011010101" => delta <= "000001111000000";
        when "00011010110" => delta <= "000001111000100";
        when "00011010111" => delta <= "000001111001000";
        when "00011011000" => delta <= "000001111001100";
        when "00011011001" => delta <= "000001111010000";
        when "00011011010" => delta <= "000001111010100";
        when "00011011011" => delta <= "000001111011000";
        when "00011011100" => delta <= "000001111011100";
        when "00011011101" => delta <= "000001111100000";
        when "00011011110" => delta <= "000001111100100";
        when "00011011111" => delta <= "000001111101001";
        when "00011100000" => delta <= "000001111101101";
        when "00011100001" => delta <= "000001111110001";
        when "00011100010" => delta <= "000001111110101";
        when "00011100011" => delta <= "000001111111001";
        when "00011100100" => delta <= "000001111111101";
        when "00011100101" => delta <= "000010000000001";
        when "00011100110" => delta <= "000010000000101";
        when "00011100111" => delta <= "000010000001001";
        when "00011101000" => delta <= "000010000001101";
        when "00011101001" => delta <= "000010000010001";
        when "00011101010" => delta <= "000010000010101";
        when "00011101011" => delta <= "000010000011001";
        when "00011101100" => delta <= "000010000011101";
        when "00011101101" => delta <= "000010000100001";
        when "00011101110" => delta <= "000010000100101";
        when "00011101111" => delta <= "000010000101001";
        when "00011110000" => delta <= "000010000101101";
        when "00011110001" => delta <= "000010000110001";
        when "00011110010" => delta <= "000010000110101";
        when "00011110011" => delta <= "000010000111000";
        when "00011110100" => delta <= "000010000111100";
        when "00011110101" => delta <= "000010001000000";
        when "00011110110" => delta <= "000010001000100";
        when "00011110111" => delta <= "000010001001000";
        when "00011111000" => delta <= "000010001001100";
        when "00011111001" => delta <= "000010001010000";
        when "00011111010" => delta <= "000010001010100";
        when "00011111011" => delta <= "000010001011000";
        when "00011111100" => delta <= "000010001011100";
        when "00011111101" => delta <= "000010001100000";
        when "00011111110" => delta <= "000010001100100";
        when "00011111111" => delta <= "000010001101000";
        when "00100000000" => delta <= "000010001101100";
        when "00100000001" => delta <= "000010001101111";
        when "00100000010" => delta <= "000010001110011";
        when "00100000011" => delta <= "000010001110111";
        when "00100000100" => delta <= "000010001111011";
        when "00100000101" => delta <= "000010001111111";
        when "00100000110" => delta <= "000010010000011";
        when "00100000111" => delta <= "000010010000111";
        when "00100001000" => delta <= "000010010001011";
        when "00100001001" => delta <= "000010010001111";
        when "00100001010" => delta <= "000010010010010";
        when "00100001011" => delta <= "000010010010110";
        when "00100001100" => delta <= "000010010011010";
        when "00100001101" => delta <= "000010010011110";
        when "00100001110" => delta <= "000010010100010";
        when "00100001111" => delta <= "000010010100110";
        when "00100010000" => delta <= "000010010101010";
        when "00100010001" => delta <= "000010010101101";
        when "00100010010" => delta <= "000010010110001";
        when "00100010011" => delta <= "000010010110101";
        when "00100010100" => delta <= "000010010111001";
        when "00100010101" => delta <= "000010010111101";
        when "00100010110" => delta <= "000010011000000";
        when "00100010111" => delta <= "000010011000100";
        when "00100011000" => delta <= "000010011001000";
        when "00100011001" => delta <= "000010011001100";
        when "00100011010" => delta <= "000010011010000";
        when "00100011011" => delta <= "000010011010011";
        when "00100011100" => delta <= "000010011010111";
        when "00100011101" => delta <= "000010011011011";
        when "00100011110" => delta <= "000010011011111";
        when "00100011111" => delta <= "000010011100011";
        when "00100100000" => delta <= "000010011100110";
        when "00100100001" => delta <= "000010011101010";
        when "00100100010" => delta <= "000010011101110";
        when "00100100011" => delta <= "000010011110010";
        when "00100100100" => delta <= "000010011110101";
        when "00100100101" => delta <= "000010011111001";
        when "00100100110" => delta <= "000010011111101";
        when "00100100111" => delta <= "000010100000001";
        when "00100101000" => delta <= "000010100000100";
        when "00100101001" => delta <= "000010100001000";
        when "00100101010" => delta <= "000010100001100";
        when "00100101011" => delta <= "000010100010000";
        when "00100101100" => delta <= "000010100010011";
        when "00100101101" => delta <= "000010100010111";
        when "00100101110" => delta <= "000010100011011";
        when "00100101111" => delta <= "000010100011111";
        when "00100110000" => delta <= "000010100100010";
        when "00100110001" => delta <= "000010100100110";
        when "00100110010" => delta <= "000010100101010";
        when "00100110011" => delta <= "000010100101101";
        when "00100110100" => delta <= "000010100110001";
        when "00100110101" => delta <= "000010100110101";
        when "00100110110" => delta <= "000010100111000";
        when "00100110111" => delta <= "000010100111100";
        when "00100111000" => delta <= "000010101000000";
        when "00100111001" => delta <= "000010101000011";
        when "00100111010" => delta <= "000010101000111";
        when "00100111011" => delta <= "000010101001011";
        when "00100111100" => delta <= "000010101001110";
        when "00100111101" => delta <= "000010101010010";
        when "00100111110" => delta <= "000010101010110";
        when "00100111111" => delta <= "000010101011001";
        when "00101000000" => delta <= "000010101011101";
        when "00101000001" => delta <= "000010101100001";
        when "00101000010" => delta <= "000010101100100";
        when "00101000011" => delta <= "000010101101000";
        when "00101000100" => delta <= "000010101101100";
        when "00101000101" => delta <= "000010101101111";
        when "00101000110" => delta <= "000010101110011";
        when "00101000111" => delta <= "000010101110110";
        when "00101001000" => delta <= "000010101111010";
        when "00101001001" => delta <= "000010101111110";
        when "00101001010" => delta <= "000010110000001";
        when "00101001011" => delta <= "000010110000101";
        when "00101001100" => delta <= "000010110001000";
        when "00101001101" => delta <= "000010110001100";
        when "00101001110" => delta <= "000010110010000";
        when "00101001111" => delta <= "000010110010011";
        when "00101010000" => delta <= "000010110010111";
        when "00101010001" => delta <= "000010110011010";
        when "00101010010" => delta <= "000010110011110";
        when "00101010011" => delta <= "000010110100001";
        when "00101010100" => delta <= "000010110100101";
        when "00101010101" => delta <= "000010110101000";
        when "00101010110" => delta <= "000010110101100";
        when "00101010111" => delta <= "000010110110000";
        when "00101011000" => delta <= "000010110110011";
        when "00101011001" => delta <= "000010110110111";
        when "00101011010" => delta <= "000010110111010";
        when "00101011011" => delta <= "000010110111110";
        when "00101011100" => delta <= "000010111000001";
        when "00101011101" => delta <= "000010111000101";
        when "00101011110" => delta <= "000010111001000";
        when "00101011111" => delta <= "000010111001100";
        when "00101100000" => delta <= "000010111001111";
        when "00101100001" => delta <= "000010111010011";
        when "00101100010" => delta <= "000010111010110";
        when "00101100011" => delta <= "000010111011010";
        when "00101100100" => delta <= "000010111011101";
        when "00101100101" => delta <= "000010111100001";
        when "00101100110" => delta <= "000010111100100";
        when "00101100111" => delta <= "000010111101000";
        when "00101101000" => delta <= "000010111101011";
        when "00101101001" => delta <= "000010111101111";
        when "00101101010" => delta <= "000010111110010";
        when "00101101011" => delta <= "000010111110110";
        when "00101101100" => delta <= "000010111111001";
        when "00101101101" => delta <= "000010111111100";
        when "00101101110" => delta <= "000011000000000";
        when "00101101111" => delta <= "000011000000011";
        when "00101110000" => delta <= "000011000000111";
        when "00101110001" => delta <= "000011000001010";
        when "00101110010" => delta <= "000011000001110";
        when "00101110011" => delta <= "000011000010001";
        when "00101110100" => delta <= "000011000010101";
        when "00101110101" => delta <= "000011000011000";
        when "00101110110" => delta <= "000011000011011";
        when "00101110111" => delta <= "000011000011111";
        when "00101111000" => delta <= "000011000100010";
        when "00101111001" => delta <= "000011000100110";
        when "00101111010" => delta <= "000011000101001";
        when "00101111011" => delta <= "000011000101100";
        when "00101111100" => delta <= "000011000110000";
        when "00101111101" => delta <= "000011000110011";
        when "00101111110" => delta <= "000011000110111";
        when "00101111111" => delta <= "000011000111010";
        when "00110000000" => delta <= "000011000111101";
        when "00110000001" => delta <= "000011001000001";
        when "00110000010" => delta <= "000011001000100";
        when "00110000011" => delta <= "000011001000111";
        when "00110000100" => delta <= "000011001001011";
        when "00110000101" => delta <= "000011001001110";
        when "00110000110" => delta <= "000011001010001";
        when "00110000111" => delta <= "000011001010101";
        when "00110001000" => delta <= "000011001011000";
        when "00110001001" => delta <= "000011001011011";
        when "00110001010" => delta <= "000011001011111";
        when "00110001011" => delta <= "000011001100010";
        when "00110001100" => delta <= "000011001100101";
        when "00110001101" => delta <= "000011001101001";
        when "00110001110" => delta <= "000011001101100";
        when "00110001111" => delta <= "000011001101111";
        when "00110010000" => delta <= "000011001110011";
        when "00110010001" => delta <= "000011001110110";
        when "00110010010" => delta <= "000011001111001";
        when "00110010011" => delta <= "000011001111100";
        when "00110010100" => delta <= "000011010000000";
        when "00110010101" => delta <= "000011010000011";
        when "00110010110" => delta <= "000011010000110";
        when "00110010111" => delta <= "000011010001010";
        when "00110011000" => delta <= "000011010001101";
        when "00110011001" => delta <= "000011010010000";
        when "00110011010" => delta <= "000011010010011";
        when "00110011011" => delta <= "000011010010111";
        when "00110011100" => delta <= "000011010011010";
        when "00110011101" => delta <= "000011010011101";
        when "00110011110" => delta <= "000011010100000";
        when "00110011111" => delta <= "000011010100100";
        when "00110100000" => delta <= "000011010100111";
        when "00110100001" => delta <= "000011010101010";
        when "00110100010" => delta <= "000011010101101";
        when "00110100011" => delta <= "000011010110001";
        when "00110100100" => delta <= "000011010110100";
        when "00110100101" => delta <= "000011010110111";
        when "00110100110" => delta <= "000011010111010";
        when "00110100111" => delta <= "000011010111101";
        when "00110101000" => delta <= "000011011000001";
        when "00110101001" => delta <= "000011011000100";
        when "00110101010" => delta <= "000011011000111";
        when "00110101011" => delta <= "000011011001010";
        when "00110101100" => delta <= "000011011001101";
        when "00110101101" => delta <= "000011011010000";
        when "00110101110" => delta <= "000011011010100";
        when "00110101111" => delta <= "000011011010111";
        when "00110110000" => delta <= "000011011011010";
        when "00110110001" => delta <= "000011011011101";
        when "00110110010" => delta <= "000011011100000";
        when "00110110011" => delta <= "000011011100011";
        when "00110110100" => delta <= "000011011100111";
        when "00110110101" => delta <= "000011011101010";
        when "00110110110" => delta <= "000011011101101";
        when "00110110111" => delta <= "000011011110000";
        when "00110111000" => delta <= "000011011110011";
        when "00110111001" => delta <= "000011011110110";
        when "00110111010" => delta <= "000011011111001";
        when "00110111011" => delta <= "000011011111100";
        when "00110111100" => delta <= "000011100000000";
        when "00110111101" => delta <= "000011100000011";
        when "00110111110" => delta <= "000011100000110";
        when "00110111111" => delta <= "000011100001001";
        when "00111000000" => delta <= "000011100001100";
        when "00111000001" => delta <= "000011100001111";
        when "00111000010" => delta <= "000011100010010";
        when "00111000011" => delta <= "000011100010101";
        when "00111000100" => delta <= "000011100011000";
        when "00111000101" => delta <= "000011100011011";
        when "00111000110" => delta <= "000011100011110";
        when "00111000111" => delta <= "000011100100010";
        when "00111001000" => delta <= "000011100100101";
        when "00111001001" => delta <= "000011100101000";
        when "00111001010" => delta <= "000011100101011";
        when "00111001011" => delta <= "000011100101110";
        when "00111001100" => delta <= "000011100110001";
        when "00111001101" => delta <= "000011100110100";
        when "00111001110" => delta <= "000011100110111";
        when "00111001111" => delta <= "000011100111010";
        when "00111010000" => delta <= "000011100111101";
        when "00111010001" => delta <= "000011101000000";
        when "00111010010" => delta <= "000011101000011";
        when "00111010011" => delta <= "000011101000110";
        when "00111010100" => delta <= "000011101001001";
        when "00111010101" => delta <= "000011101001100";
        when "00111010110" => delta <= "000011101001111";
        when "00111010111" => delta <= "000011101010010";
        when "00111011000" => delta <= "000011101010101";
        when "00111011001" => delta <= "000011101011000";
        when "00111011010" => delta <= "000011101011011";
        when "00111011011" => delta <= "000011101011110";
        when "00111011100" => delta <= "000011101100001";
        when "00111011101" => delta <= "000011101100100";
        when "00111011110" => delta <= "000011101100111";
        when "00111011111" => delta <= "000011101101010";
        when "00111100000" => delta <= "000011101101101";
        when "00111100001" => delta <= "000011101110000";
        when "00111100010" => delta <= "000011101110011";
        when "00111100011" => delta <= "000011101110110";
        when "00111100100" => delta <= "000011101111000";
        when "00111100101" => delta <= "000011101111011";
        when "00111100110" => delta <= "000011101111110";
        when "00111100111" => delta <= "000011110000001";
        when "00111101000" => delta <= "000011110000100";
        when "00111101001" => delta <= "000011110000111";
        when "00111101010" => delta <= "000011110001010";
        when "00111101011" => delta <= "000011110001101";
        when "00111101100" => delta <= "000011110010000";
        when "00111101101" => delta <= "000011110010011";
        when "00111101110" => delta <= "000011110010110";
        when "00111101111" => delta <= "000011110011000";
        when "00111110000" => delta <= "000011110011011";
        when "00111110001" => delta <= "000011110011110";
        when "00111110010" => delta <= "000011110100001";
        when "00111110011" => delta <= "000011110100100";
        when "00111110100" => delta <= "000011110100111";
        when "00111110101" => delta <= "000011110101010";
        when "00111110110" => delta <= "000011110101101";
        when "00111110111" => delta <= "000011110101111";
        when "00111111000" => delta <= "000011110110010";
        when "00111111001" => delta <= "000011110110101";
        when "00111111010" => delta <= "000011110111000";
        when "00111111011" => delta <= "000011110111011";
        when "00111111100" => delta <= "000011110111110";
        when "00111111101" => delta <= "000011111000000";
        when "00111111110" => delta <= "000011111000011";
        when "00111111111" => delta <= "000011111000110";
        when "01000000000" => delta <= "000011111001001";
        when "01000000001" => delta <= "000011111001100";
        when "01000000010" => delta <= "000011111001110";
        when "01000000011" => delta <= "000011111010001";
        when "01000000100" => delta <= "000011111010100";
        when "01000000101" => delta <= "000011111010111";
        when "01000000110" => delta <= "000011111011010";
        when "01000000111" => delta <= "000011111011100";
        when "01000001000" => delta <= "000011111011111";
        when "01000001001" => delta <= "000011111100010";
        when "01000001010" => delta <= "000011111100101";
        when "01000001011" => delta <= "000011111101000";
        when "01000001100" => delta <= "000011111101010";
        when "01000001101" => delta <= "000011111101101";
        when "01000001110" => delta <= "000011111110000";
        when "01000001111" => delta <= "000011111110011";
        when "01000010000" => delta <= "000011111110101";
        when "01000010001" => delta <= "000011111111000";
        when "01000010010" => delta <= "000011111111011";
        when "01000010011" => delta <= "000011111111101";
        when "01000010100" => delta <= "000100000000000";
        when "01000010101" => delta <= "000100000000011";
        when "01000010110" => delta <= "000100000000110";
        when "01000010111" => delta <= "000100000001000";
        when "01000011000" => delta <= "000100000001011";
        when "01000011001" => delta <= "000100000001110";
        when "01000011010" => delta <= "000100000010000";
        when "01000011011" => delta <= "000100000010011";
        when "01000011100" => delta <= "000100000010110";
        when "01000011101" => delta <= "000100000011000";
        when "01000011110" => delta <= "000100000011011";
        when "01000011111" => delta <= "000100000011110";
        when "01000100000" => delta <= "000100000100000";
        when "01000100001" => delta <= "000100000100011";
        when "01000100010" => delta <= "000100000100110";
        when "01000100011" => delta <= "000100000101000";
        when "01000100100" => delta <= "000100000101011";
        when "01000100101" => delta <= "000100000101110";
        when "01000100110" => delta <= "000100000110000";
        when "01000100111" => delta <= "000100000110011";
        when "01000101000" => delta <= "000100000110110";
        when "01000101001" => delta <= "000100000111000";
        when "01000101010" => delta <= "000100000111011";
        when "01000101011" => delta <= "000100000111110";
        when "01000101100" => delta <= "000100001000000";
        when "01000101101" => delta <= "000100001000011";
        when "01000101110" => delta <= "000100001000101";
        when "01000101111" => delta <= "000100001001000";
        when "01000110000" => delta <= "000100001001011";
        when "01000110001" => delta <= "000100001001101";
        when "01000110010" => delta <= "000100001010000";
        when "01000110011" => delta <= "000100001010010";
        when "01000110100" => delta <= "000100001010101";
        when "01000110101" => delta <= "000100001010111";
        when "01000110110" => delta <= "000100001011010";
        when "01000110111" => delta <= "000100001011101";
        when "01000111000" => delta <= "000100001011111";
        when "01000111001" => delta <= "000100001100010";
        when "01000111010" => delta <= "000100001100100";
        when "01000111011" => delta <= "000100001100111";
        when "01000111100" => delta <= "000100001101001";
        when "01000111101" => delta <= "000100001101100";
        when "01000111110" => delta <= "000100001101110";
        when "01000111111" => delta <= "000100001110001";
        when "01001000000" => delta <= "000100001110011";
        when "01001000001" => delta <= "000100001110110";
        when "01001000010" => delta <= "000100001111000";
        when "01001000011" => delta <= "000100001111011";
        when "01001000100" => delta <= "000100001111110";
        when "01001000101" => delta <= "000100010000000";
        when "01001000110" => delta <= "000100010000010";
        when "01001000111" => delta <= "000100010000101";
        when "01001001000" => delta <= "000100010000111";
        when "01001001001" => delta <= "000100010001010";
        when "01001001010" => delta <= "000100010001100";
        when "01001001011" => delta <= "000100010001111";
        when "01001001100" => delta <= "000100010010001";
        when "01001001101" => delta <= "000100010010100";
        when "01001001110" => delta <= "000100010010110";
        when "01001001111" => delta <= "000100010011001";
        when "01001010000" => delta <= "000100010011011";
        when "01001010001" => delta <= "000100010011110";
        when "01001010010" => delta <= "000100010100000";
        when "01001010011" => delta <= "000100010100011";
        when "01001010100" => delta <= "000100010100101";
        when "01001010101" => delta <= "000100010100111";
        when "01001010110" => delta <= "000100010101010";
        when "01001010111" => delta <= "000100010101100";
        when "01001011000" => delta <= "000100010101111";
        when "01001011001" => delta <= "000100010110001";
        when "01001011010" => delta <= "000100010110011";
        when "01001011011" => delta <= "000100010110110";
        when "01001011100" => delta <= "000100010111000";
        when "01001011101" => delta <= "000100010111011";
        when "01001011110" => delta <= "000100010111101";
        when "01001011111" => delta <= "000100010111111";
        when "01001100000" => delta <= "000100011000010";
        when "01001100001" => delta <= "000100011000100";
        when "01001100010" => delta <= "000100011000111";
        when "01001100011" => delta <= "000100011001001";
        when "01001100100" => delta <= "000100011001011";
        when "01001100101" => delta <= "000100011001110";
        when "01001100110" => delta <= "000100011010000";
        when "01001100111" => delta <= "000100011010010";
        when "01001101000" => delta <= "000100011010101";
        when "01001101001" => delta <= "000100011010111";
        when "01001101010" => delta <= "000100011011001";
        when "01001101011" => delta <= "000100011011100";
        when "01001101100" => delta <= "000100011011110";
        when "01001101101" => delta <= "000100011100000";
        when "01001101110" => delta <= "000100011100011";
        when "01001101111" => delta <= "000100011100101";
        when "01001110000" => delta <= "000100011100111";
        when "01001110001" => delta <= "000100011101001";
        when "01001110010" => delta <= "000100011101100";
        when "01001110011" => delta <= "000100011101110";
        when "01001110100" => delta <= "000100011110000";
        when "01001110101" => delta <= "000100011110011";
        when "01001110110" => delta <= "000100011110101";
        when "01001110111" => delta <= "000100011110111";
        when "01001111000" => delta <= "000100011111001";
        when "01001111001" => delta <= "000100011111100";
        when "01001111010" => delta <= "000100011111110";
        when "01001111011" => delta <= "000100100000000";
        when "01001111100" => delta <= "000100100000010";
        when "01001111101" => delta <= "000100100000101";
        when "01001111110" => delta <= "000100100000111";
        when "01001111111" => delta <= "000100100001001";
        when "01010000000" => delta <= "000100100001011";
        when "01010000001" => delta <= "000100100001110";
        when "01010000010" => delta <= "000100100010000";
        when "01010000011" => delta <= "000100100010010";
        when "01010000100" => delta <= "000100100010100";
        when "01010000101" => delta <= "000100100010110";
        when "01010000110" => delta <= "000100100011001";
        when "01010000111" => delta <= "000100100011011";
        when "01010001000" => delta <= "000100100011101";
        when "01010001001" => delta <= "000100100011111";
        when "01010001010" => delta <= "000100100100001";
        when "01010001011" => delta <= "000100100100100";
        when "01010001100" => delta <= "000100100100110";
        when "01010001101" => delta <= "000100100101000";
        when "01010001110" => delta <= "000100100101010";
        when "01010001111" => delta <= "000100100101100";
        when "01010010000" => delta <= "000100100101110";
        when "01010010001" => delta <= "000100100110000";
        when "01010010010" => delta <= "000100100110011";
        when "01010010011" => delta <= "000100100110101";
        when "01010010100" => delta <= "000100100110111";
        when "01010010101" => delta <= "000100100111001";
        when "01010010110" => delta <= "000100100111011";
        when "01010010111" => delta <= "000100100111101";
        when "01010011000" => delta <= "000100100111111";
        when "01010011001" => delta <= "000100101000010";
        when "01010011010" => delta <= "000100101000100";
        when "01010011011" => delta <= "000100101000110";
        when "01010011100" => delta <= "000100101001000";
        when "01010011101" => delta <= "000100101001010";
        when "01010011110" => delta <= "000100101001100";
        when "01010011111" => delta <= "000100101001110";
        when "01010100000" => delta <= "000100101010000";
        when "01010100001" => delta <= "000100101010010";
        when "01010100010" => delta <= "000100101010100";
        when "01010100011" => delta <= "000100101010110";
        when "01010100100" => delta <= "000100101011000";
        when "01010100101" => delta <= "000100101011010";
        when "01010100110" => delta <= "000100101011101";
        when "01010100111" => delta <= "000100101011111";
        when "01010101000" => delta <= "000100101100001";
        when "01010101001" => delta <= "000100101100011";
        when "01010101010" => delta <= "000100101100101";
        when "01010101011" => delta <= "000100101100111";
        when "01010101100" => delta <= "000100101101001";
        when "01010101101" => delta <= "000100101101011";
        when "01010101110" => delta <= "000100101101101";
        when "01010101111" => delta <= "000100101101111";
        when "01010110000" => delta <= "000100101110001";
        when "01010110001" => delta <= "000100101110011";
        when "01010110010" => delta <= "000100101110101";
        when "01010110011" => delta <= "000100101110111";
        when "01010110100" => delta <= "000100101111001";
        when "01010110101" => delta <= "000100101111011";
        when "01010110110" => delta <= "000100101111101";
        when "01010110111" => delta <= "000100101111111";
        when "01010111000" => delta <= "000100110000001";
        when "01010111001" => delta <= "000100110000011";
        when "01010111010" => delta <= "000100110000101";
        when "01010111011" => delta <= "000100110000110";
        when "01010111100" => delta <= "000100110001000";
        when "01010111101" => delta <= "000100110001010";
        when "01010111110" => delta <= "000100110001100";
        when "01010111111" => delta <= "000100110001110";
        when "01011000000" => delta <= "000100110010000";
        when "01011000001" => delta <= "000100110010010";
        when "01011000010" => delta <= "000100110010100";
        when "01011000011" => delta <= "000100110010110";
        when "01011000100" => delta <= "000100110011000";
        when "01011000101" => delta <= "000100110011010";
        when "01011000110" => delta <= "000100110011100";
        when "01011000111" => delta <= "000100110011101";
        when "01011001000" => delta <= "000100110011111";
        when "01011001001" => delta <= "000100110100001";
        when "01011001010" => delta <= "000100110100011";
        when "01011001011" => delta <= "000100110100101";
        when "01011001100" => delta <= "000100110100111";
        when "01011001101" => delta <= "000100110101001";
        when "01011001110" => delta <= "000100110101011";
        when "01011001111" => delta <= "000100110101100";
        when "01011010000" => delta <= "000100110101110";
        when "01011010001" => delta <= "000100110110000";
        when "01011010010" => delta <= "000100110110010";
        when "01011010011" => delta <= "000100110110100";
        when "01011010100" => delta <= "000100110110110";
        when "01011010101" => delta <= "000100110110111";
        when "01011010110" => delta <= "000100110111001";
        when "01011010111" => delta <= "000100110111011";
        when "01011011000" => delta <= "000100110111101";
        when "01011011001" => delta <= "000100110111111";
        when "01011011010" => delta <= "000100111000001";
        when "01011011011" => delta <= "000100111000010";
        when "01011011100" => delta <= "000100111000100";
        when "01011011101" => delta <= "000100111000110";
        when "01011011110" => delta <= "000100111001000";
        when "01011011111" => delta <= "000100111001001";
        when "01011100000" => delta <= "000100111001011";
        when "01011100001" => delta <= "000100111001101";
        when "01011100010" => delta <= "000100111001111";
        when "01011100011" => delta <= "000100111010001";
        when "01011100100" => delta <= "000100111010010";
        when "01011100101" => delta <= "000100111010100";
        when "01011100110" => delta <= "000100111010110";
        when "01011100111" => delta <= "000100111011000";
        when "01011101000" => delta <= "000100111011001";
        when "01011101001" => delta <= "000100111011011";
        when "01011101010" => delta <= "000100111011101";
        when "01011101011" => delta <= "000100111011110";
        when "01011101100" => delta <= "000100111100000";
        when "01011101101" => delta <= "000100111100010";
        when "01011101110" => delta <= "000100111100100";
        when "01011101111" => delta <= "000100111100101";
        when "01011110000" => delta <= "000100111100111";
        when "01011110001" => delta <= "000100111101001";
        when "01011110010" => delta <= "000100111101010";
        when "01011110011" => delta <= "000100111101100";
        when "01011110100" => delta <= "000100111101110";
        when "01011110101" => delta <= "000100111101111";
        when "01011110110" => delta <= "000100111110001";
        when "01011110111" => delta <= "000100111110011";
        when "01011111000" => delta <= "000100111110100";
        when "01011111001" => delta <= "000100111110110";
        when "01011111010" => delta <= "000100111111000";
        when "01011111011" => delta <= "000100111111001";
        when "01011111100" => delta <= "000100111111011";
        when "01011111101" => delta <= "000100111111101";
        when "01011111110" => delta <= "000100111111110";
        when "01011111111" => delta <= "000101000000000";
        when "01100000000" => delta <= "000101000000001";
        when "01100000001" => delta <= "000101000000011";
        when "01100000010" => delta <= "000101000000101";
        when "01100000011" => delta <= "000101000000110";
        when "01100000100" => delta <= "000101000001000";
        when "01100000101" => delta <= "000101000001001";
        when "01100000110" => delta <= "000101000001011";
        when "01100000111" => delta <= "000101000001101";
        when "01100001000" => delta <= "000101000001110";
        when "01100001001" => delta <= "000101000010000";
        when "01100001010" => delta <= "000101000010001";
        when "01100001011" => delta <= "000101000010011";
        when "01100001100" => delta <= "000101000010100";
        when "01100001101" => delta <= "000101000010110";
        when "01100001110" => delta <= "000101000011000";
        when "01100001111" => delta <= "000101000011001";
        when "01100010000" => delta <= "000101000011011";
        when "01100010001" => delta <= "000101000011100";
        when "01100010010" => delta <= "000101000011110";
        when "01100010011" => delta <= "000101000011111";
        when "01100010100" => delta <= "000101000100001";
        when "01100010101" => delta <= "000101000100010";
        when "01100010110" => delta <= "000101000100100";
        when "01100010111" => delta <= "000101000100101";
        when "01100011000" => delta <= "000101000100111";
        when "01100011001" => delta <= "000101000101000";
        when "01100011010" => delta <= "000101000101010";
        when "01100011011" => delta <= "000101000101011";
        when "01100011100" => delta <= "000101000101101";
        when "01100011101" => delta <= "000101000101110";
        when "01100011110" => delta <= "000101000110000";
        when "01100011111" => delta <= "000101000110001";
        when "01100100000" => delta <= "000101000110011";
        when "01100100001" => delta <= "000101000110100";
        when "01100100010" => delta <= "000101000110110";
        when "01100100011" => delta <= "000101000110111";
        when "01100100100" => delta <= "000101000111000";
        when "01100100101" => delta <= "000101000111010";
        when "01100100110" => delta <= "000101000111011";
        when "01100100111" => delta <= "000101000111101";
        when "01100101000" => delta <= "000101000111110";
        when "01100101001" => delta <= "000101001000000";
        when "01100101010" => delta <= "000101001000001";
        when "01100101011" => delta <= "000101001000010";
        when "01100101100" => delta <= "000101001000100";
        when "01100101101" => delta <= "000101001000101";
        when "01100101110" => delta <= "000101001000111";
        when "01100101111" => delta <= "000101001001000";
        when "01100110000" => delta <= "000101001001001";
        when "01100110001" => delta <= "000101001001011";
        when "01100110010" => delta <= "000101001001100";
        when "01100110011" => delta <= "000101001001101";
        when "01100110100" => delta <= "000101001001111";
        when "01100110101" => delta <= "000101001010000";
        when "01100110110" => delta <= "000101001010010";
        when "01100110111" => delta <= "000101001010011";
        when "01100111000" => delta <= "000101001010100";
        when "01100111001" => delta <= "000101001010110";
        when "01100111010" => delta <= "000101001010111";
        when "01100111011" => delta <= "000101001011000";
        when "01100111100" => delta <= "000101001011010";
        when "01100111101" => delta <= "000101001011011";
        when "01100111110" => delta <= "000101001011100";
        when "01100111111" => delta <= "000101001011101";
        when "01101000000" => delta <= "000101001011111";
        when "01101000001" => delta <= "000101001100000";
        when "01101000010" => delta <= "000101001100001";
        when "01101000011" => delta <= "000101001100011";
        when "01101000100" => delta <= "000101001100100";
        when "01101000101" => delta <= "000101001100101";
        when "01101000110" => delta <= "000101001100110";
        when "01101000111" => delta <= "000101001101000";
        when "01101001000" => delta <= "000101001101001";
        when "01101001001" => delta <= "000101001101010";
        when "01101001010" => delta <= "000101001101100";
        when "01101001011" => delta <= "000101001101101";
        when "01101001100" => delta <= "000101001101110";
        when "01101001101" => delta <= "000101001101111";
        when "01101001110" => delta <= "000101001110000";
        when "01101001111" => delta <= "000101001110010";
        when "01101010000" => delta <= "000101001110011";
        when "01101010001" => delta <= "000101001110100";
        when "01101010010" => delta <= "000101001110101";
        when "01101010011" => delta <= "000101001110111";
        when "01101010100" => delta <= "000101001111000";
        when "01101010101" => delta <= "000101001111001";
        when "01101010110" => delta <= "000101001111010";
        when "01101010111" => delta <= "000101001111011";
        when "01101011000" => delta <= "000101001111101";
        when "01101011001" => delta <= "000101001111110";
        when "01101011010" => delta <= "000101001111111";
        when "01101011011" => delta <= "000101010000000";
        when "01101011100" => delta <= "000101010000001";
        when "01101011101" => delta <= "000101010000010";
        when "01101011110" => delta <= "000101010000100";
        when "01101011111" => delta <= "000101010000101";
        when "01101100000" => delta <= "000101010000110";
        when "01101100001" => delta <= "000101010000111";
        when "01101100010" => delta <= "000101010001000";
        when "01101100011" => delta <= "000101010001001";
        when "01101100100" => delta <= "000101010001010";
        when "01101100101" => delta <= "000101010001011";
        when "01101100110" => delta <= "000101010001101";
        when "01101100111" => delta <= "000101010001110";
        when "01101101000" => delta <= "000101010001111";
        when "01101101001" => delta <= "000101010010000";
        when "01101101010" => delta <= "000101010010001";
        when "01101101011" => delta <= "000101010010010";
        when "01101101100" => delta <= "000101010010011";
        when "01101101101" => delta <= "000101010010100";
        when "01101101110" => delta <= "000101010010101";
        when "01101101111" => delta <= "000101010010110";
        when "01101110000" => delta <= "000101010010111";
        when "01101110001" => delta <= "000101010011000";
        when "01101110010" => delta <= "000101010011010";
        when "01101110011" => delta <= "000101010011011";
        when "01101110100" => delta <= "000101010011100";
        when "01101110101" => delta <= "000101010011101";
        when "01101110110" => delta <= "000101010011110";
        when "01101110111" => delta <= "000101010011111";
        when "01101111000" => delta <= "000101010100000";
        when "01101111001" => delta <= "000101010100001";
        when "01101111010" => delta <= "000101010100010";
        when "01101111011" => delta <= "000101010100011";
        when "01101111100" => delta <= "000101010100100";
        when "01101111101" => delta <= "000101010100101";
        when "01101111110" => delta <= "000101010100110";
        when "01101111111" => delta <= "000101010100111";
        when "01110000000" => delta <= "000101010101000";
        when "01110000001" => delta <= "000101010101001";
        when "01110000010" => delta <= "000101010101010";
        when "01110000011" => delta <= "000101010101011";
        when "01110000100" => delta <= "000101010101100";
        when "01110000101" => delta <= "000101010101101";
        when "01110000110" => delta <= "000101010101101";
        when "01110000111" => delta <= "000101010101110";
        when "01110001000" => delta <= "000101010101111";
        when "01110001001" => delta <= "000101010110000";
        when "01110001010" => delta <= "000101010110001";
        when "01110001011" => delta <= "000101010110010";
        when "01110001100" => delta <= "000101010110011";
        when "01110001101" => delta <= "000101010110100";
        when "01110001110" => delta <= "000101010110101";
        when "01110001111" => delta <= "000101010110110";
        when "01110010000" => delta <= "000101010110111";
        when "01110010001" => delta <= "000101010111000";
        when "01110010010" => delta <= "000101010111000";
        when "01110010011" => delta <= "000101010111001";
        when "01110010100" => delta <= "000101010111010";
        when "01110010101" => delta <= "000101010111011";
        when "01110010110" => delta <= "000101010111100";
        when "01110010111" => delta <= "000101010111101";
        when "01110011000" => delta <= "000101010111110";
        when "01110011001" => delta <= "000101010111111";
        when "01110011010" => delta <= "000101010111111";
        when "01110011011" => delta <= "000101011000000";
        when "01110011100" => delta <= "000101011000001";
        when "01110011101" => delta <= "000101011000010";
        when "01110011110" => delta <= "000101011000011";
        when "01110011111" => delta <= "000101011000100";
        when "01110100000" => delta <= "000101011000100";
        when "01110100001" => delta <= "000101011000101";
        when "01110100010" => delta <= "000101011000110";
        when "01110100011" => delta <= "000101011000111";
        when "01110100100" => delta <= "000101011001000";
        when "01110100101" => delta <= "000101011001000";
        when "01110100110" => delta <= "000101011001001";
        when "01110100111" => delta <= "000101011001010";
        when "01110101000" => delta <= "000101011001011";
        when "01110101001" => delta <= "000101011001100";
        when "01110101010" => delta <= "000101011001100";
        when "01110101011" => delta <= "000101011001101";
        when "01110101100" => delta <= "000101011001110";
        when "01110101101" => delta <= "000101011001111";
        when "01110101110" => delta <= "000101011001111";
        when "01110101111" => delta <= "000101011010000";
        when "01110110000" => delta <= "000101011010001";
        when "01110110001" => delta <= "000101011010010";
        when "01110110010" => delta <= "000101011010010";
        when "01110110011" => delta <= "000101011010011";
        when "01110110100" => delta <= "000101011010100";
        when "01110110101" => delta <= "000101011010100";
        when "01110110110" => delta <= "000101011010101";
        when "01110110111" => delta <= "000101011010110";
        when "01110111000" => delta <= "000101011010110";
        when "01110111001" => delta <= "000101011010111";
        when "01110111010" => delta <= "000101011011000";
        when "01110111011" => delta <= "000101011011001";
        when "01110111100" => delta <= "000101011011001";
        when "01110111101" => delta <= "000101011011010";
        when "01110111110" => delta <= "000101011011011";
        when "01110111111" => delta <= "000101011011011";
        when "01111000000" => delta <= "000101011011100";
        when "01111000001" => delta <= "000101011011100";
        when "01111000010" => delta <= "000101011011101";
        when "01111000011" => delta <= "000101011011110";
        when "01111000100" => delta <= "000101011011110";
        when "01111000101" => delta <= "000101011011111";
        when "01111000110" => delta <= "000101011100000";
        when "01111000111" => delta <= "000101011100000";
        when "01111001000" => delta <= "000101011100001";
        when "01111001001" => delta <= "000101011100001";
        when "01111001010" => delta <= "000101011100010";
        when "01111001011" => delta <= "000101011100011";
        when "01111001100" => delta <= "000101011100011";
        when "01111001101" => delta <= "000101011100100";
        when "01111001110" => delta <= "000101011100100";
        when "01111001111" => delta <= "000101011100101";
        when "01111010000" => delta <= "000101011100110";
        when "01111010001" => delta <= "000101011100110";
        when "01111010010" => delta <= "000101011100111";
        when "01111010011" => delta <= "000101011100111";
        when "01111010100" => delta <= "000101011101000";
        when "01111010101" => delta <= "000101011101000";
        when "01111010110" => delta <= "000101011101001";
        when "01111010111" => delta <= "000101011101001";
        when "01111011000" => delta <= "000101011101010";
        when "01111011001" => delta <= "000101011101010";
        when "01111011010" => delta <= "000101011101011";
        when "01111011011" => delta <= "000101011101011";
        when "01111011100" => delta <= "000101011101100";
        when "01111011101" => delta <= "000101011101100";
        when "01111011110" => delta <= "000101011101101";
        when "01111011111" => delta <= "000101011101101";
        when "01111100000" => delta <= "000101011101110";
        when "01111100001" => delta <= "000101011101110";
        when "01111100010" => delta <= "000101011101111";
        when "01111100011" => delta <= "000101011101111";
        when "01111100100" => delta <= "000101011110000";
        when "01111100101" => delta <= "000101011110000";
        when "01111100110" => delta <= "000101011110001";
        when "01111100111" => delta <= "000101011110001";
        when "01111101000" => delta <= "000101011110010";
        when "01111101001" => delta <= "000101011110010";
        when "01111101010" => delta <= "000101011110011";
        when "01111101011" => delta <= "000101011110011";
        when "01111101100" => delta <= "000101011110011";
        when "01111101101" => delta <= "000101011110100";
        when "01111101110" => delta <= "000101011110100";
        when "01111101111" => delta <= "000101011110101";
        when "01111110000" => delta <= "000101011110101";
        when "01111110001" => delta <= "000101011110101";
        when "01111110010" => delta <= "000101011110110";
        when "01111110011" => delta <= "000101011110110";
        when "01111110100" => delta <= "000101011110111";
        when "01111110101" => delta <= "000101011110111";
        when "01111110110" => delta <= "000101011110111";
        when "01111110111" => delta <= "000101011111000";
        when "01111111000" => delta <= "000101011111000";
        when "01111111001" => delta <= "000101011111000";
        when "01111111010" => delta <= "000101011111001";
        when "01111111011" => delta <= "000101011111001";
        when "01111111100" => delta <= "000101011111001";
        when "01111111101" => delta <= "000101011111010";
        when "01111111110" => delta <= "000101011111010";
        when "01111111111" => delta <= "000101011111010";
        when "10000000000" => delta <= "000101011111011";
        when "10000000001" => delta <= "000101011111011";
        when "10000000010" => delta <= "000101011111011";
        when "10000000011" => delta <= "000101011111100";
        when "10000000100" => delta <= "000101011111100";
        when "10000000101" => delta <= "000101011111100";
        when "10000000110" => delta <= "000101011111100";
        when "10000000111" => delta <= "000101011111101";
        when "10000001000" => delta <= "000101011111101";
        when "10000001001" => delta <= "000101011111101";
        when "10000001010" => delta <= "000101011111110";
        when "10000001011" => delta <= "000101011111110";
        when "10000001100" => delta <= "000101011111110";
        when "10000001101" => delta <= "000101011111110";
        when "10000001110" => delta <= "000101011111111";
        when "10000001111" => delta <= "000101011111111";
        when "10000010000" => delta <= "000101011111111";
        when "10000010001" => delta <= "000101011111111";
        when "10000010010" => delta <= "000101011111111";
        when "10000010011" => delta <= "000101100000000";
        when "10000010100" => delta <= "000101100000000";
        when "10000010101" => delta <= "000101100000000";
        when "10000010110" => delta <= "000101100000000";
        when "10000010111" => delta <= "000101100000000";
        when "10000011000" => delta <= "000101100000001";
        when "10000011001" => delta <= "000101100000001";
        when "10000011010" => delta <= "000101100000001";
        when "10000011011" => delta <= "000101100000001";
        when "10000011100" => delta <= "000101100000001";
        when "10000011101" => delta <= "000101100000010";
        when "10000011110" => delta <= "000101100000010";
        when "10000011111" => delta <= "000101100000010";
        when "10000100000" => delta <= "000101100000010";
        when "10000100001" => delta <= "000101100000010";
        when "10000100010" => delta <= "000101100000010";
        when "10000100011" => delta <= "000101100000010";
        when "10000100100" => delta <= "000101100000011";
        when "10000100101" => delta <= "000101100000011";
        when "10000100110" => delta <= "000101100000011";
        when "10000100111" => delta <= "000101100000011";
        when "10000101000" => delta <= "000101100000011";
        when "10000101001" => delta <= "000101100000011";
        when "10000101010" => delta <= "000101100000011";
        when "10000101011" => delta <= "000101100000011";
        when "10000101100" => delta <= "000101100000011";
        when "10000101101" => delta <= "000101100000011";
        when "10000101110" => delta <= "000101100000011";
        when "10000101111" => delta <= "000101100000100";
        when "10000110000" => delta <= "000101100000100";
        when "10000110001" => delta <= "000101100000100";
        when "10000110010" => delta <= "000101100000100";
        when "10000110011" => delta <= "000101100000100";
        when "10000110100" => delta <= "000101100000100";
        when "10000110101" => delta <= "000101100000100";
        when "10000110110" => delta <= "000101100000100";
        when "10000110111" => delta <= "000101100000100";
        when "10000111000" => delta <= "000101100000100";
        when "10000111001" => delta <= "000101100000100";
        when "10000111010" => delta <= "000101100000100";
        when "10000111011" => delta <= "000101100000100";
        when "10000111100" => delta <= "000101100000100";
        when "10000111101" => delta <= "000101100000100";
        when "10000111110" => delta <= "000101100000100";
        when "10000111111" => delta <= "000101100000100";
        when "10001000000" => delta <= "000101100000100";
        when "10001000001" => delta <= "000101100000100";
        when "10001000010" => delta <= "000101100000100";
        when "10001000011" => delta <= "000101100000100";
        when "10001000100" => delta <= "000101100000100";
        when "10001000101" => delta <= "000101100000100";
        when "10001000110" => delta <= "000101100000100";
        when "10001000111" => delta <= "000101100000011";
        when "10001001000" => delta <= "000101100000011";
        when "10001001001" => delta <= "000101100000011";
        when "10001001010" => delta <= "000101100000011";
        when "10001001011" => delta <= "000101100000011";
        when "10001001100" => delta <= "000101100000011";
        when "10001001101" => delta <= "000101100000011";
        when "10001001110" => delta <= "000101100000011";
        when "10001001111" => delta <= "000101100000011";
        when "10001010000" => delta <= "000101100000011";
        when "10001010001" => delta <= "000101100000011";
        when "10001010010" => delta <= "000101100000010";
        when "10001010011" => delta <= "000101100000010";
        when "10001010100" => delta <= "000101100000010";
        when "10001010101" => delta <= "000101100000010";
        when "10001010110" => delta <= "000101100000010";
        when "10001010111" => delta <= "000101100000010";
        when "10001011000" => delta <= "000101100000010";
        when "10001011001" => delta <= "000101100000001";
        when "10001011010" => delta <= "000101100000001";
        when "10001011011" => delta <= "000101100000001";
        when "10001011100" => delta <= "000101100000001";
        when "10001011101" => delta <= "000101100000001";
        when "10001011110" => delta <= "000101100000000";
        when "10001011111" => delta <= "000101100000000";
        when "10001100000" => delta <= "000101100000000";
        when "10001100001" => delta <= "000101100000000";
        when "10001100010" => delta <= "000101100000000";
        when "10001100011" => delta <= "000101011111111";
        when "10001100100" => delta <= "000101011111111";
        when "10001100101" => delta <= "000101011111111";
        when "10001100110" => delta <= "000101011111111";
        when "10001100111" => delta <= "000101011111110";
        when "10001101000" => delta <= "000101011111110";
        when "10001101001" => delta <= "000101011111110";
        when "10001101010" => delta <= "000101011111110";
        when "10001101011" => delta <= "000101011111101";
        when "10001101100" => delta <= "000101011111101";
        when "10001101101" => delta <= "000101011111101";
        when "10001101110" => delta <= "000101011111101";
        when "10001101111" => delta <= "000101011111100";
        when "10001110000" => delta <= "000101011111100";
        when "10001110001" => delta <= "000101011111100";
        when "10001110010" => delta <= "000101011111011";
        when "10001110011" => delta <= "000101011111011";
        when "10001110100" => delta <= "000101011111011";
        when "10001110101" => delta <= "000101011111011";
        when "10001110110" => delta <= "000101011111010";
        when "10001110111" => delta <= "000101011111010";
        when "10001111000" => delta <= "000101011111010";
        when "10001111001" => delta <= "000101011111001";
        when "10001111010" => delta <= "000101011111001";
        when "10001111011" => delta <= "000101011111001";
        when "10001111100" => delta <= "000101011111000";
        when "10001111101" => delta <= "000101011111000";
        when "10001111110" => delta <= "000101011110111";
        when "10001111111" => delta <= "000101011110111";
        when "10010000000" => delta <= "000101011110111";
        when "10010000001" => delta <= "000101011110110";
        when "10010000010" => delta <= "000101011110110";
        when "10010000011" => delta <= "000101011110110";
        when "10010000100" => delta <= "000101011110101";
        when "10010000101" => delta <= "000101011110101";
        when "10010000110" => delta <= "000101011110100";
        when "10010000111" => delta <= "000101011110100";
        when "10010001000" => delta <= "000101011110011";
        when "10010001001" => delta <= "000101011110011";
        when "10010001010" => delta <= "000101011110011";
        when "10010001011" => delta <= "000101011110010";
        when "10010001100" => delta <= "000101011110010";
        when "10010001101" => delta <= "000101011110001";
        when "10010001110" => delta <= "000101011110001";
        when "10010001111" => delta <= "000101011110000";
        when "10010010000" => delta <= "000101011110000";
        when "10010010001" => delta <= "000101011101111";
        when "10010010010" => delta <= "000101011101111";
        when "10010010011" => delta <= "000101011101110";
        when "10010010100" => delta <= "000101011101110";
        when "10010010101" => delta <= "000101011101101";
        when "10010010110" => delta <= "000101011101101";
        when "10010010111" => delta <= "000101011101100";
        when "10010011000" => delta <= "000101011101100";
        when "10010011001" => delta <= "000101011101011";
        when "10010011010" => delta <= "000101011101011";
        when "10010011011" => delta <= "000101011101010";
        when "10010011100" => delta <= "000101011101010";
        when "10010011101" => delta <= "000101011101001";
        when "10010011110" => delta <= "000101011101001";
        when "10010011111" => delta <= "000101011101000";
        when "10010100000" => delta <= "000101011101000";
        when "10010100001" => delta <= "000101011100111";
        when "10010100010" => delta <= "000101011100111";
        when "10010100011" => delta <= "000101011100110";
        when "10010100100" => delta <= "000101011100101";
        when "10010100101" => delta <= "000101011100101";
        when "10010100110" => delta <= "000101011100100";
        when "10010100111" => delta <= "000101011100100";
        when "10010101000" => delta <= "000101011100011";
        when "10010101001" => delta <= "000101011100010";
        when "10010101010" => delta <= "000101011100010";
        when "10010101011" => delta <= "000101011100001";
        when "10010101100" => delta <= "000101011100001";
        when "10010101101" => delta <= "000101011100000";
        when "10010101110" => delta <= "000101011011111";
        when "10010101111" => delta <= "000101011011111";
        when "10010110000" => delta <= "000101011011110";
        when "10010110001" => delta <= "000101011011101";
        when "10010110010" => delta <= "000101011011101";
        when "10010110011" => delta <= "000101011011100";
        when "10010110100" => delta <= "000101011011011";
        when "10010110101" => delta <= "000101011011011";
        when "10010110110" => delta <= "000101011011010";
        when "10010110111" => delta <= "000101011011001";
        when "10010111000" => delta <= "000101011011001";
        when "10010111001" => delta <= "000101011011000";
        when "10010111010" => delta <= "000101011010111";
        when "10010111011" => delta <= "000101011010110";
        when "10010111100" => delta <= "000101011010110";
        when "10010111101" => delta <= "000101011010101";
        when "10010111110" => delta <= "000101011010100";
        when "10010111111" => delta <= "000101011010100";
        when "10011000000" => delta <= "000101011010011";
        when "10011000001" => delta <= "000101011010010";
        when "10011000010" => delta <= "000101011010001";
        when "10011000011" => delta <= "000101011010001";
        when "10011000100" => delta <= "000101011010000";
        when "10011000101" => delta <= "000101011001111";
        when "10011000110" => delta <= "000101011001110";
        when "10011000111" => delta <= "000101011001110";
        when "10011001000" => delta <= "000101011001101";
        when "10011001001" => delta <= "000101011001100";
        when "10011001010" => delta <= "000101011001011";
        when "10011001011" => delta <= "000101011001010";
        when "10011001100" => delta <= "000101011001010";
        when "10011001101" => delta <= "000101011001001";
        when "10011001110" => delta <= "000101011001000";
        when "10011001111" => delta <= "000101011000111";
        when "10011010000" => delta <= "000101011000110";
        when "10011010001" => delta <= "000101011000101";
        when "10011010010" => delta <= "000101011000101";
        when "10011010011" => delta <= "000101011000100";
        when "10011010100" => delta <= "000101011000011";
        when "10011010101" => delta <= "000101011000010";
        when "10011010110" => delta <= "000101011000001";
        when "10011010111" => delta <= "000101011000000";
        when "10011011000" => delta <= "000101010111111";
        when "10011011001" => delta <= "000101010111111";
        when "10011011010" => delta <= "000101010111110";
        when "10011011011" => delta <= "000101010111101";
        when "10011011100" => delta <= "000101010111100";
        when "10011011101" => delta <= "000101010111011";
        when "10011011110" => delta <= "000101010111010";
        when "10011011111" => delta <= "000101010111001";
        when "10011100000" => delta <= "000101010111000";
        when "10011100001" => delta <= "000101010110111";
        when "10011100010" => delta <= "000101010110110";
        when "10011100011" => delta <= "000101010110101";
        when "10011100100" => delta <= "000101010110101";
        when "10011100101" => delta <= "000101010110100";
        when "10011100110" => delta <= "000101010110011";
        when "10011100111" => delta <= "000101010110010";
        when "10011101000" => delta <= "000101010110001";
        when "10011101001" => delta <= "000101010110000";
        when "10011101010" => delta <= "000101010101111";
        when "10011101011" => delta <= "000101010101110";
        when "10011101100" => delta <= "000101010101101";
        when "10011101101" => delta <= "000101010101100";
        when "10011101110" => delta <= "000101010101011";
        when "10011101111" => delta <= "000101010101010";
        when "10011110000" => delta <= "000101010101001";
        when "10011110001" => delta <= "000101010101000";
        when "10011110010" => delta <= "000101010100111";
        when "10011110011" => delta <= "000101010100110";
        when "10011110100" => delta <= "000101010100101";
        when "10011110101" => delta <= "000101010100100";
        when "10011110110" => delta <= "000101010100011";
        when "10011110111" => delta <= "000101010100010";
        when "10011111000" => delta <= "000101010100000";
        when "10011111001" => delta <= "000101010011111";
        when "10011111010" => delta <= "000101010011110";
        when "10011111011" => delta <= "000101010011101";
        when "10011111100" => delta <= "000101010011100";
        when "10011111101" => delta <= "000101010011011";
        when "10011111110" => delta <= "000101010011010";
        when "10011111111" => delta <= "000101010011001";
        when "10100000000" => delta <= "000101010011000";
        when "10100000001" => delta <= "000101010010111";
        when "10100000010" => delta <= "000101010010110";
        when "10100000011" => delta <= "000101010010100";
        when "10100000100" => delta <= "000101010010011";
        when "10100000101" => delta <= "000101010010010";
        when "10100000110" => delta <= "000101010010001";
        when "10100000111" => delta <= "000101010010000";
        when "10100001000" => delta <= "000101010001111";
        when "10100001001" => delta <= "000101010001110";
        when "10100001010" => delta <= "000101010001100";
        when "10100001011" => delta <= "000101010001011";
        when "10100001100" => delta <= "000101010001010";
        when "10100001101" => delta <= "000101010001001";
        when "10100001110" => delta <= "000101010001000";
        when "10100001111" => delta <= "000101010000111";
        when "10100010000" => delta <= "000101010000101";
        when "10100010001" => delta <= "000101010000100";
        when "10100010010" => delta <= "000101010000011";
        when "10100010011" => delta <= "000101010000010";
        when "10100010100" => delta <= "000101010000001";
        when "10100010101" => delta <= "000101001111111";
        when "10100010110" => delta <= "000101001111110";
        when "10100010111" => delta <= "000101001111101";
        when "10100011000" => delta <= "000101001111100";
        when "10100011001" => delta <= "000101001111010";
        when "10100011010" => delta <= "000101001111001";
        when "10100011011" => delta <= "000101001111000";
        when "10100011100" => delta <= "000101001110111";
        when "10100011101" => delta <= "000101001110101";
        when "10100011110" => delta <= "000101001110100";
        when "10100011111" => delta <= "000101001110011";
        when "10100100000" => delta <= "000101001110001";
        when "10100100001" => delta <= "000101001110000";
        when "10100100010" => delta <= "000101001101111";
        when "10100100011" => delta <= "000101001101110";
        when "10100100100" => delta <= "000101001101100";
        when "10100100101" => delta <= "000101001101011";
        when "10100100110" => delta <= "000101001101010";
        when "10100100111" => delta <= "000101001101000";
        when "10100101000" => delta <= "000101001100111";
        when "10100101001" => delta <= "000101001100110";
        when "10100101010" => delta <= "000101001100100";
        when "10100101011" => delta <= "000101001100011";
        when "10100101100" => delta <= "000101001100010";
        when "10100101101" => delta <= "000101001100000";
        when "10100101110" => delta <= "000101001011111";
        when "10100101111" => delta <= "000101001011101";
        when "10100110000" => delta <= "000101001011100";
        when "10100110001" => delta <= "000101001011011";
        when "10100110010" => delta <= "000101001011001";
        when "10100110011" => delta <= "000101001011000";
        when "10100110100" => delta <= "000101001010110";
        when "10100110101" => delta <= "000101001010101";
        when "10100110110" => delta <= "000101001010100";
        when "10100110111" => delta <= "000101001010010";
        when "10100111000" => delta <= "000101001010001";
        when "10100111001" => delta <= "000101001001111";
        when "10100111010" => delta <= "000101001001110";
        when "10100111011" => delta <= "000101001001100";
        when "10100111100" => delta <= "000101001001011";
        when "10100111101" => delta <= "000101001001001";
        when "10100111110" => delta <= "000101001001000";
        when "10100111111" => delta <= "000101001000111";
        when "10101000000" => delta <= "000101001000101";
        when "10101000001" => delta <= "000101001000100";
        when "10101000010" => delta <= "000101001000010";
        when "10101000011" => delta <= "000101001000001";
        when "10101000100" => delta <= "000101000111111";
        when "10101000101" => delta <= "000101000111110";
        when "10101000110" => delta <= "000101000111100";
        when "10101000111" => delta <= "000101000111011";
        when "10101001000" => delta <= "000101000111001";
        when "10101001001" => delta <= "000101000110111";
        when "10101001010" => delta <= "000101000110110";
        when "10101001011" => delta <= "000101000110100";
        when "10101001100" => delta <= "000101000110011";
        when "10101001101" => delta <= "000101000110001";
        when "10101001110" => delta <= "000101000110000";
        when "10101001111" => delta <= "000101000101110";
        when "10101010000" => delta <= "000101000101101";
        when "10101010001" => delta <= "000101000101011";
        when "10101010010" => delta <= "000101000101001";
        when "10101010011" => delta <= "000101000101000";
        when "10101010100" => delta <= "000101000100110";
        when "10101010101" => delta <= "000101000100101";
        when "10101010110" => delta <= "000101000100011";
        when "10101010111" => delta <= "000101000100001";
        when "10101011000" => delta <= "000101000100000";
        when "10101011001" => delta <= "000101000011110";
        when "10101011010" => delta <= "000101000011101";
        when "10101011011" => delta <= "000101000011011";
        when "10101011100" => delta <= "000101000011001";
        when "10101011101" => delta <= "000101000011000";
        when "10101011110" => delta <= "000101000010110";
        when "10101011111" => delta <= "000101000010100";
        when "10101100000" => delta <= "000101000010011";
        when "10101100001" => delta <= "000101000010001";
        when "10101100010" => delta <= "000101000001111";
        when "10101100011" => delta <= "000101000001110";
        when "10101100100" => delta <= "000101000001100";
        when "10101100101" => delta <= "000101000001010";
        when "10101100110" => delta <= "000101000001000";
        when "10101100111" => delta <= "000101000000111";
        when "10101101000" => delta <= "000101000000101";
        when "10101101001" => delta <= "000101000000011";
        when "10101101010" => delta <= "000101000000010";
        when "10101101011" => delta <= "000101000000000";
        when "10101101100" => delta <= "000100111111110";
        when "10101101101" => delta <= "000100111111100";
        when "10101101110" => delta <= "000100111111011";
        when "10101101111" => delta <= "000100111111001";
        when "10101110000" => delta <= "000100111110111";
        when "10101110001" => delta <= "000100111110101";
        when "10101110010" => delta <= "000100111110100";
        when "10101110011" => delta <= "000100111110010";
        when "10101110100" => delta <= "000100111110000";
        when "10101110101" => delta <= "000100111101110";
        when "10101110110" => delta <= "000100111101100";
        when "10101110111" => delta <= "000100111101011";
        when "10101111000" => delta <= "000100111101001";
        when "10101111001" => delta <= "000100111100111";
        when "10101111010" => delta <= "000100111100101";
        when "10101111011" => delta <= "000100111100011";
        when "10101111100" => delta <= "000100111100001";
        when "10101111101" => delta <= "000100111100000";
        when "10101111110" => delta <= "000100111011110";
        when "10101111111" => delta <= "000100111011100";
        when "10110000000" => delta <= "000100111011010";
        when "10110000001" => delta <= "000100111011000";
        when "10110000010" => delta <= "000100111010110";
        when "10110000011" => delta <= "000100111010100";
        when "10110000100" => delta <= "000100111010011";
        when "10110000101" => delta <= "000100111010001";
        when "10110000110" => delta <= "000100111001111";
        when "10110000111" => delta <= "000100111001101";
        when "10110001000" => delta <= "000100111001011";
        when "10110001001" => delta <= "000100111001001";
        when "10110001010" => delta <= "000100111000111";
        when "10110001011" => delta <= "000100111000101";
        when "10110001100" => delta <= "000100111000011";
        when "10110001101" => delta <= "000100111000001";
        when "10110001110" => delta <= "000100110111111";
        when "10110001111" => delta <= "000100110111101";
        when "10110010000" => delta <= "000100110111011";
        when "10110010001" => delta <= "000100110111010";
        when "10110010010" => delta <= "000100110111000";
        when "10110010011" => delta <= "000100110110110";
        when "10110010100" => delta <= "000100110110100";
        when "10110010101" => delta <= "000100110110010";
        when "10110010110" => delta <= "000100110110000";
        when "10110010111" => delta <= "000100110101110";
        when "10110011000" => delta <= "000100110101100";
        when "10110011001" => delta <= "000100110101010";
        when "10110011010" => delta <= "000100110101000";
        when "10110011011" => delta <= "000100110100110";
        when "10110011100" => delta <= "000100110100100";
        when "10110011101" => delta <= "000100110100001";
        when "10110011110" => delta <= "000100110011111";
        when "10110011111" => delta <= "000100110011101";
        when "10110100000" => delta <= "000100110011011";
        when "10110100001" => delta <= "000100110011001";
        when "10110100010" => delta <= "000100110010111";
        when "10110100011" => delta <= "000100110010101";
        when "10110100100" => delta <= "000100110010011";
        when "10110100101" => delta <= "000100110010001";
        when "10110100110" => delta <= "000100110001111";
        when "10110100111" => delta <= "000100110001101";
        when "10110101000" => delta <= "000100110001011";
        when "10110101001" => delta <= "000100110001001";
        when "10110101010" => delta <= "000100110000110";
        when "10110101011" => delta <= "000100110000100";
        when "10110101100" => delta <= "000100110000010";
        when "10110101101" => delta <= "000100110000000";
        when "10110101110" => delta <= "000100101111110";
        when "10110101111" => delta <= "000100101111100";
        when "10110110000" => delta <= "000100101111010";
        when "10110110001" => delta <= "000100101110111";
        when "10110110010" => delta <= "000100101110101";
        when "10110110011" => delta <= "000100101110011";
        when "10110110100" => delta <= "000100101110001";
        when "10110110101" => delta <= "000100101101111";
        when "10110110110" => delta <= "000100101101101";
        when "10110110111" => delta <= "000100101101010";
        when "10110111000" => delta <= "000100101101000";
        when "10110111001" => delta <= "000100101100110";
        when "10110111010" => delta <= "000100101100100";
        when "10110111011" => delta <= "000100101100010";
        when "10110111100" => delta <= "000100101011111";
        when "10110111101" => delta <= "000100101011101";
        when "10110111110" => delta <= "000100101011011";
        when "10110111111" => delta <= "000100101011001";
        when "10111000000" => delta <= "000100101010110";
        when "10111000001" => delta <= "000100101010100";
        when "10111000010" => delta <= "000100101010010";
        when "10111000011" => delta <= "000100101010000";
        when "10111000100" => delta <= "000100101001101";
        when "10111000101" => delta <= "000100101001011";
        when "10111000110" => delta <= "000100101001001";
        when "10111000111" => delta <= "000100101000110";
        when "10111001000" => delta <= "000100101000100";
        when "10111001001" => delta <= "000100101000010";
        when "10111001010" => delta <= "000100100111111";
        when "10111001011" => delta <= "000100100111101";
        when "10111001100" => delta <= "000100100111011";
        when "10111001101" => delta <= "000100100111000";
        when "10111001110" => delta <= "000100100110110";
        when "10111001111" => delta <= "000100100110100";
        when "10111010000" => delta <= "000100100110001";
        when "10111010001" => delta <= "000100100101111";
        when "10111010010" => delta <= "000100100101101";
        when "10111010011" => delta <= "000100100101010";
        when "10111010100" => delta <= "000100100101000";
        when "10111010101" => delta <= "000100100100110";
        when "10111010110" => delta <= "000100100100011";
        when "10111010111" => delta <= "000100100100001";
        when "10111011000" => delta <= "000100100011110";
        when "10111011001" => delta <= "000100100011100";
        when "10111011010" => delta <= "000100100011010";
        when "10111011011" => delta <= "000100100010111";
        when "10111011100" => delta <= "000100100010101";
        when "10111011101" => delta <= "000100100010010";
        when "10111011110" => delta <= "000100100010000";
        when "10111011111" => delta <= "000100100001101";
        when "10111100000" => delta <= "000100100001011";
        when "10111100001" => delta <= "000100100001001";
        when "10111100010" => delta <= "000100100000110";
        when "10111100011" => delta <= "000100100000100";
        when "10111100100" => delta <= "000100100000001";
        when "10111100101" => delta <= "000100011111111";
        when "10111100110" => delta <= "000100011111100";
        when "10111100111" => delta <= "000100011111010";
        when "10111101000" => delta <= "000100011110111";
        when "10111101001" => delta <= "000100011110101";
        when "10111101010" => delta <= "000100011110010";
        when "10111101011" => delta <= "000100011110000";
        when "10111101100" => delta <= "000100011101101";
        when "10111101101" => delta <= "000100011101011";
        when "10111101110" => delta <= "000100011101000";
        when "10111101111" => delta <= "000100011100101";
        when "10111110000" => delta <= "000100011100011";
        when "10111110001" => delta <= "000100011100000";
        when "10111110010" => delta <= "000100011011110";
        when "10111110011" => delta <= "000100011011011";
        when "10111110100" => delta <= "000100011011001";
        when "10111110101" => delta <= "000100011010110";
        when "10111110110" => delta <= "000100011010011";
        when "10111110111" => delta <= "000100011010001";
        when "10111111000" => delta <= "000100011001110";
        when "10111111001" => delta <= "000100011001100";
        when "10111111010" => delta <= "000100011001001";
        when "10111111011" => delta <= "000100011000110";
        when "10111111100" => delta <= "000100011000100";
        when "10111111101" => delta <= "000100011000001";
        when "10111111110" => delta <= "000100010111111";
        when "10111111111" => delta <= "000100010111100";
        when "11000000000" => delta <= "000100010111001";
        when "11000000001" => delta <= "000100010110111";
        when "11000000010" => delta <= "000100010110100";
        when "11000000011" => delta <= "000100010110001";
        when "11000000100" => delta <= "000100010101111";
        when "11000000101" => delta <= "000100010101100";
        when "11000000110" => delta <= "000100010101001";
        when "11000000111" => delta <= "000100010100111";
        when "11000001000" => delta <= "000100010100100";
        when "11000001001" => delta <= "000100010100001";
        when "11000001010" => delta <= "000100010011110";
        when "11000001011" => delta <= "000100010011100";
        when "11000001100" => delta <= "000100010011001";
        when "11000001101" => delta <= "000100010010110";
        when "11000001110" => delta <= "000100010010011";
        when "11000001111" => delta <= "000100010010001";
        when "11000010000" => delta <= "000100010001110";
        when "11000010001" => delta <= "000100010001011";
        when "11000010010" => delta <= "000100010001000";
        when "11000010011" => delta <= "000100010000110";
        when "11000010100" => delta <= "000100010000011";
        when "11000010101" => delta <= "000100010000000";
        when "11000010110" => delta <= "000100001111101";
        when "11000010111" => delta <= "000100001111011";
        when "11000011000" => delta <= "000100001111000";
        when "11000011001" => delta <= "000100001110101";
        when "11000011010" => delta <= "000100001110010";
        when "11000011011" => delta <= "000100001101111";
        when "11000011100" => delta <= "000100001101100";
        when "11000011101" => delta <= "000100001101010";
        when "11000011110" => delta <= "000100001100111";
        when "11000011111" => delta <= "000100001100100";
        when "11000100000" => delta <= "000100001100001";
        when "11000100001" => delta <= "000100001011110";
        when "11000100010" => delta <= "000100001011011";
        when "11000100011" => delta <= "000100001011000";
        when "11000100100" => delta <= "000100001010110";
        when "11000100101" => delta <= "000100001010011";
        when "11000100110" => delta <= "000100001010000";
        when "11000100111" => delta <= "000100001001101";
        when "11000101000" => delta <= "000100001001010";
        when "11000101001" => delta <= "000100001000111";
        when "11000101010" => delta <= "000100001000100";
        when "11000101011" => delta <= "000100001000001";
        when "11000101100" => delta <= "000100000111110";
        when "11000101101" => delta <= "000100000111011";
        when "11000101110" => delta <= "000100000111000";
        when "11000101111" => delta <= "000100000110101";
        when "11000110000" => delta <= "000100000110011";
        when "11000110001" => delta <= "000100000110000";
        when "11000110010" => delta <= "000100000101101";
        when "11000110011" => delta <= "000100000101010";
        when "11000110100" => delta <= "000100000100111";
        when "11000110101" => delta <= "000100000100100";
        when "11000110110" => delta <= "000100000100001";
        when "11000110111" => delta <= "000100000011110";
        when "11000111000" => delta <= "000100000011011";
        when "11000111001" => delta <= "000100000011000";
        when "11000111010" => delta <= "000100000010101";
        when "11000111011" => delta <= "000100000010010";
        when "11000111100" => delta <= "000100000001111";
        when "11000111101" => delta <= "000100000001100";
        when "11000111110" => delta <= "000100000001000";
        when "11000111111" => delta <= "000100000000101";
        when "11001000000" => delta <= "000100000000010";
        when "11001000001" => delta <= "000011111111111";
        when "11001000010" => delta <= "000011111111100";
        when "11001000011" => delta <= "000011111111001";
        when "11001000100" => delta <= "000011111110110";
        when "11001000101" => delta <= "000011111110011";
        when "11001000110" => delta <= "000011111110000";
        when "11001000111" => delta <= "000011111101101";
        when "11001001000" => delta <= "000011111101010";
        when "11001001001" => delta <= "000011111100111";
        when "11001001010" => delta <= "000011111100011";
        when "11001001011" => delta <= "000011111100000";
        when "11001001100" => delta <= "000011111011101";
        when "11001001101" => delta <= "000011111011010";
        when "11001001110" => delta <= "000011111010111";
        when "11001001111" => delta <= "000011111010100";
        when "11001010000" => delta <= "000011111010001";
        when "11001010001" => delta <= "000011111001101";
        when "11001010010" => delta <= "000011111001010";
        when "11001010011" => delta <= "000011111000111";
        when "11001010100" => delta <= "000011111000100";
        when "11001010101" => delta <= "000011111000001";
        when "11001010110" => delta <= "000011110111101";
        when "11001010111" => delta <= "000011110111010";
        when "11001011000" => delta <= "000011110110111";
        when "11001011001" => delta <= "000011110110100";
        when "11001011010" => delta <= "000011110110001";
        when "11001011011" => delta <= "000011110101101";
        when "11001011100" => delta <= "000011110101010";
        when "11001011101" => delta <= "000011110100111";
        when "11001011110" => delta <= "000011110100100";
        when "11001011111" => delta <= "000011110100000";
        when "11001100000" => delta <= "000011110011101";
        when "11001100001" => delta <= "000011110011010";
        when "11001100010" => delta <= "000011110010110";
        when "11001100011" => delta <= "000011110010011";
        when "11001100100" => delta <= "000011110010000";
        when "11001100101" => delta <= "000011110001101";
        when "11001100110" => delta <= "000011110001001";
        when "11001100111" => delta <= "000011110000110";
        when "11001101000" => delta <= "000011110000011";
        when "11001101001" => delta <= "000011101111111";
        when "11001101010" => delta <= "000011101111100";
        when "11001101011" => delta <= "000011101111001";
        when "11001101100" => delta <= "000011101110101";
        when "11001101101" => delta <= "000011101110010";
        when "11001101110" => delta <= "000011101101111";
        when "11001101111" => delta <= "000011101101011";
        when "11001110000" => delta <= "000011101101000";
        when "11001110001" => delta <= "000011101100100";
        when "11001110010" => delta <= "000011101100001";
        when "11001110011" => delta <= "000011101011110";
        when "11001110100" => delta <= "000011101011010";
        when "11001110101" => delta <= "000011101010111";
        when "11001110110" => delta <= "000011101010011";
        when "11001110111" => delta <= "000011101010000";
        when "11001111000" => delta <= "000011101001101";
        when "11001111001" => delta <= "000011101001001";
        when "11001111010" => delta <= "000011101000110";
        when "11001111011" => delta <= "000011101000010";
        when "11001111100" => delta <= "000011100111111";
        when "11001111101" => delta <= "000011100111011";
        when "11001111110" => delta <= "000011100111000";
        when "11001111111" => delta <= "000011100110100";
        when "11010000000" => delta <= "000011100110001";
        when "11010000001" => delta <= "000011100101110";
        when "11010000010" => delta <= "000011100101010";
        when "11010000011" => delta <= "000011100100111";
        when "11010000100" => delta <= "000011100100011";
        when "11010000101" => delta <= "000011100100000";
        when "11010000110" => delta <= "000011100011100";
        when "11010000111" => delta <= "000011100011000";
        when "11010001000" => delta <= "000011100010101";
        when "11010001001" => delta <= "000011100010001";
        when "11010001010" => delta <= "000011100001110";
        when "11010001011" => delta <= "000011100001010";
        when "11010001100" => delta <= "000011100000111";
        when "11010001101" => delta <= "000011100000011";
        when "11010001110" => delta <= "000011100000000";
        when "11010001111" => delta <= "000011011111100";
        when "11010010000" => delta <= "000011011111000";
        when "11010010001" => delta <= "000011011110101";
        when "11010010010" => delta <= "000011011110001";
        when "11010010011" => delta <= "000011011101110";
        when "11010010100" => delta <= "000011011101010";
        when "11010010101" => delta <= "000011011100110";
        when "11010010110" => delta <= "000011011100011";
        when "11010010111" => delta <= "000011011011111";
        when "11010011000" => delta <= "000011011011100";
        when "11010011001" => delta <= "000011011011000";
        when "11010011010" => delta <= "000011011010100";
        when "11010011011" => delta <= "000011011010001";
        when "11010011100" => delta <= "000011011001101";
        when "11010011101" => delta <= "000011011001001";
        when "11010011110" => delta <= "000011011000110";
        when "11010011111" => delta <= "000011011000010";
        when "11010100000" => delta <= "000011010111110";
        when "11010100001" => delta <= "000011010111011";
        when "11010100010" => delta <= "000011010110111";
        when "11010100011" => delta <= "000011010110011";
        when "11010100100" => delta <= "000011010101111";
        when "11010100101" => delta <= "000011010101100";
        when "11010100110" => delta <= "000011010101000";
        when "11010100111" => delta <= "000011010100100";
        when "11010101000" => delta <= "000011010100000";
        when "11010101001" => delta <= "000011010011101";
        when "11010101010" => delta <= "000011010011001";
        when "11010101011" => delta <= "000011010010101";
        when "11010101100" => delta <= "000011010010001";
        when "11010101101" => delta <= "000011010001110";
        when "11010101110" => delta <= "000011010001010";
        when "11010101111" => delta <= "000011010000110";
        when "11010110000" => delta <= "000011010000010";
        when "11010110001" => delta <= "000011001111110";
        when "11010110010" => delta <= "000011001111011";
        when "11010110011" => delta <= "000011001110111";
        when "11010110100" => delta <= "000011001110011";
        when "11010110101" => delta <= "000011001101111";
        when "11010110110" => delta <= "000011001101011";
        when "11010110111" => delta <= "000011001101000";
        when "11010111000" => delta <= "000011001100100";
        when "11010111001" => delta <= "000011001100000";
        when "11010111010" => delta <= "000011001011100";
        when "11010111011" => delta <= "000011001011000";
        when "11010111100" => delta <= "000011001010100";
        when "11010111101" => delta <= "000011001010000";
        when "11010111110" => delta <= "000011001001100";
        when "11010111111" => delta <= "000011001001001";
        when "11011000000" => delta <= "000011001000101";
        when "11011000001" => delta <= "000011001000001";
        when "11011000010" => delta <= "000011000111101";
        when "11011000011" => delta <= "000011000111001";
        when "11011000100" => delta <= "000011000110101";
        when "11011000101" => delta <= "000011000110001";
        when "11011000110" => delta <= "000011000101101";
        when "11011000111" => delta <= "000011000101001";
        when "11011001000" => delta <= "000011000100101";
        when "11011001001" => delta <= "000011000100001";
        when "11011001010" => delta <= "000011000011101";
        when "11011001011" => delta <= "000011000011001";
        when "11011001100" => delta <= "000011000010101";
        when "11011001101" => delta <= "000011000010001";
        when "11011001110" => delta <= "000011000001101";
        when "11011001111" => delta <= "000011000001001";
        when "11011010000" => delta <= "000011000000101";
        when "11011010001" => delta <= "000011000000001";
        when "11011010010" => delta <= "000010111111101";
        when "11011010011" => delta <= "000010111111001";
        when "11011010100" => delta <= "000010111110101";
        when "11011010101" => delta <= "000010111110001";
        when "11011010110" => delta <= "000010111101101";
        when "11011010111" => delta <= "000010111101001";
        when "11011011000" => delta <= "000010111100101";
        when "11011011001" => delta <= "000010111100001";
        when "11011011010" => delta <= "000010111011101";
        when "11011011011" => delta <= "000010111011001";
        when "11011011100" => delta <= "000010111010101";
        when "11011011101" => delta <= "000010111010000";
        when "11011011110" => delta <= "000010111001100";
        when "11011011111" => delta <= "000010111001000";
        when "11011100000" => delta <= "000010111000100";
        when "11011100001" => delta <= "000010111000000";
        when "11011100010" => delta <= "000010110111100";
        when "11011100011" => delta <= "000010110111000";
        when "11011100100" => delta <= "000010110110100";
        when "11011100101" => delta <= "000010110101111";
        when "11011100110" => delta <= "000010110101011";
        when "11011100111" => delta <= "000010110100111";
        when "11011101000" => delta <= "000010110100011";
        when "11011101001" => delta <= "000010110011111";
        when "11011101010" => delta <= "000010110011011";
        when "11011101011" => delta <= "000010110010110";
        when "11011101100" => delta <= "000010110010010";
        when "11011101101" => delta <= "000010110001110";
        when "11011101110" => delta <= "000010110001010";
        when "11011101111" => delta <= "000010110000110";
        when "11011110000" => delta <= "000010110000001";
        when "11011110001" => delta <= "000010101111101";
        when "11011110010" => delta <= "000010101111001";
        when "11011110011" => delta <= "000010101110101";
        when "11011110100" => delta <= "000010101110000";
        when "11011110101" => delta <= "000010101101100";
        when "11011110110" => delta <= "000010101101000";
        when "11011110111" => delta <= "000010101100011";
        when "11011111000" => delta <= "000010101011111";
        when "11011111001" => delta <= "000010101011011";
        when "11011111010" => delta <= "000010101010111";
        when "11011111011" => delta <= "000010101010010";
        when "11011111100" => delta <= "000010101001110";
        when "11011111101" => delta <= "000010101001010";
        when "11011111110" => delta <= "000010101000101";
        when "11011111111" => delta <= "000010101000001";
        when "11100000000" => delta <= "000010100111101";
        when "11100000001" => delta <= "000010100111000";
        when "11100000010" => delta <= "000010100110100";
        when "11100000011" => delta <= "000010100110000";
        when "11100000100" => delta <= "000010100101011";
        when "11100000101" => delta <= "000010100100111";
        when "11100000110" => delta <= "000010100100011";
        when "11100000111" => delta <= "000010100011110";
        when "11100001000" => delta <= "000010100011010";
        when "11100001001" => delta <= "000010100010101";
        when "11100001010" => delta <= "000010100010001";
        when "11100001011" => delta <= "000010100001100";
        when "11100001100" => delta <= "000010100001000";
        when "11100001101" => delta <= "000010100000100";
        when "11100001110" => delta <= "000010011111111";
        when "11100001111" => delta <= "000010011111011";
        when "11100010000" => delta <= "000010011110110";
        when "11100010001" => delta <= "000010011110010";
        when "11100010010" => delta <= "000010011101101";
        when "11100010011" => delta <= "000010011101001";
        when "11100010100" => delta <= "000010011100100";
        when "11100010101" => delta <= "000010011100000";
        when "11100010110" => delta <= "000010011011011";
        when "11100010111" => delta <= "000010011010111";
        when "11100011000" => delta <= "000010011010010";
        when "11100011001" => delta <= "000010011001110";
        when "11100011010" => delta <= "000010011001001";
        when "11100011011" => delta <= "000010011000101";
        when "11100011100" => delta <= "000010011000000";
        when "11100011101" => delta <= "000010010111100";
        when "11100011110" => delta <= "000010010110111";
        when "11100011111" => delta <= "000010010110011";
        when "11100100000" => delta <= "000010010101110";
        when "11100100001" => delta <= "000010010101010";
        when "11100100010" => delta <= "000010010100101";
        when "11100100011" => delta <= "000010010100000";
        when "11100100100" => delta <= "000010010011100";
        when "11100100101" => delta <= "000010010010111";
        when "11100100110" => delta <= "000010010010011";
        when "11100100111" => delta <= "000010010001110";
        when "11100101000" => delta <= "000010010001001";
        when "11100101001" => delta <= "000010010000101";
        when "11100101010" => delta <= "000010010000000";
        when "11100101011" => delta <= "000010001111100";
        when "11100101100" => delta <= "000010001110111";
        when "11100101101" => delta <= "000010001110010";
        when "11100101110" => delta <= "000010001101110";
        when "11100101111" => delta <= "000010001101001";
        when "11100110000" => delta <= "000010001100100";
        when "11100110001" => delta <= "000010001100000";
        when "11100110010" => delta <= "000010001011011";
        when "11100110011" => delta <= "000010001010110";
        when "11100110100" => delta <= "000010001010001";
        when "11100110101" => delta <= "000010001001101";
        when "11100110110" => delta <= "000010001001000";
        when "11100110111" => delta <= "000010001000011";
        when "11100111000" => delta <= "000010000111111";
        when "11100111001" => delta <= "000010000111010";
        when "11100111010" => delta <= "000010000110101";
        when "11100111011" => delta <= "000010000110000";
        when "11100111100" => delta <= "000010000101100";
        when "11100111101" => delta <= "000010000100111";
        when "11100111110" => delta <= "000010000100010";
        when "11100111111" => delta <= "000010000011101";
        when "11101000000" => delta <= "000010000011001";
        when "11101000001" => delta <= "000010000010100";
        when "11101000010" => delta <= "000010000001111";
        when "11101000011" => delta <= "000010000001010";
        when "11101000100" => delta <= "000010000000101";
        when "11101000101" => delta <= "000010000000001";
        when "11101000110" => delta <= "000001111111100";
        when "11101000111" => delta <= "000001111110111";
        when "11101001000" => delta <= "000001111110010";
        when "11101001001" => delta <= "000001111101101";
        when "11101001010" => delta <= "000001111101000";
        when "11101001011" => delta <= "000001111100011";
        when "11101001100" => delta <= "000001111011111";
        when "11101001101" => delta <= "000001111011010";
        when "11101001110" => delta <= "000001111010101";
        when "11101001111" => delta <= "000001111010000";
        when "11101010000" => delta <= "000001111001011";
        when "11101010001" => delta <= "000001111000110";
        when "11101010010" => delta <= "000001111000001";
        when "11101010011" => delta <= "000001110111100";
        when "11101010100" => delta <= "000001110110111";
        when "11101010101" => delta <= "000001110110010";
        when "11101010110" => delta <= "000001110101101";
        when "11101010111" => delta <= "000001110101001";
        when "11101011000" => delta <= "000001110100100";
        when "11101011001" => delta <= "000001110011111";
        when "11101011010" => delta <= "000001110011010";
        when "11101011011" => delta <= "000001110010101";
        when "11101011100" => delta <= "000001110010000";
        when "11101011101" => delta <= "000001110001011";
        when "11101011110" => delta <= "000001110000110";
        when "11101011111" => delta <= "000001110000001";
        when "11101100000" => delta <= "000001101111100";
        when "11101100001" => delta <= "000001101110111";
        when "11101100010" => delta <= "000001101110010";
        when "11101100011" => delta <= "000001101101101";
        when "11101100100" => delta <= "000001101101000";
        when "11101100101" => delta <= "000001101100011";
        when "11101100110" => delta <= "000001101011101";
        when "11101100111" => delta <= "000001101011000";
        when "11101101000" => delta <= "000001101010011";
        when "11101101001" => delta <= "000001101001110";
        when "11101101010" => delta <= "000001101001001";
        when "11101101011" => delta <= "000001101000100";
        when "11101101100" => delta <= "000001100111111";
        when "11101101101" => delta <= "000001100111010";
        when "11101101110" => delta <= "000001100110101";
        when "11101101111" => delta <= "000001100110000";
        when "11101110000" => delta <= "000001100101011";
        when "11101110001" => delta <= "000001100100101";
        when "11101110010" => delta <= "000001100100000";
        when "11101110011" => delta <= "000001100011011";
        when "11101110100" => delta <= "000001100010110";
        when "11101110101" => delta <= "000001100010001";
        when "11101110110" => delta <= "000001100001100";
        when "11101110111" => delta <= "000001100000110";
        when "11101111000" => delta <= "000001100000001";
        when "11101111001" => delta <= "000001011111100";
        when "11101111010" => delta <= "000001011110111";
        when "11101111011" => delta <= "000001011110010";
        when "11101111100" => delta <= "000001011101100";
        when "11101111101" => delta <= "000001011100111";
        when "11101111110" => delta <= "000001011100010";
        when "11101111111" => delta <= "000001011011101";
        when "11110000000" => delta <= "000001011011000";
        when "11110000001" => delta <= "000001011010010";
        when "11110000010" => delta <= "000001011001101";
        when "11110000011" => delta <= "000001011001000";
        when "11110000100" => delta <= "000001011000011";
        when "11110000101" => delta <= "000001010111101";
        when "11110000110" => delta <= "000001010111000";
        when "11110000111" => delta <= "000001010110011";
        when "11110001000" => delta <= "000001010101101";
        when "11110001001" => delta <= "000001010101000";
        when "11110001010" => delta <= "000001010100011";
        when "11110001011" => delta <= "000001010011101";
        when "11110001100" => delta <= "000001010011000";
        when "11110001101" => delta <= "000001010010011";
        when "11110001110" => delta <= "000001010001101";
        when "11110001111" => delta <= "000001010001000";
        when "11110010000" => delta <= "000001010000011";
        when "11110010001" => delta <= "000001001111101";
        when "11110010010" => delta <= "000001001111000";
        when "11110010011" => delta <= "000001001110011";
        when "11110010100" => delta <= "000001001101101";
        when "11110010101" => delta <= "000001001101000";
        when "11110010110" => delta <= "000001001100010";
        when "11110010111" => delta <= "000001001011101";
        when "11110011000" => delta <= "000001001011000";
        when "11110011001" => delta <= "000001001010010";
        when "11110011010" => delta <= "000001001001101";
        when "11110011011" => delta <= "000001001000111";
        when "11110011100" => delta <= "000001001000010";
        when "11110011101" => delta <= "000001000111100";
        when "11110011110" => delta <= "000001000110111";
        when "11110011111" => delta <= "000001000110010";
        when "11110100000" => delta <= "000001000101100";
        when "11110100001" => delta <= "000001000100111";
        when "11110100010" => delta <= "000001000100001";
        when "11110100011" => delta <= "000001000011100";
        when "11110100100" => delta <= "000001000010110";
        when "11110100101" => delta <= "000001000010001";
        when "11110100110" => delta <= "000001000001011";
        when "11110100111" => delta <= "000001000000110";
        when "11110101000" => delta <= "000001000000000";
        when "11110101001" => delta <= "000000111111010";
        when "11110101010" => delta <= "000000111110101";
        when "11110101011" => delta <= "000000111101111";
        when "11110101100" => delta <= "000000111101010";
        when "11110101101" => delta <= "000000111100100";
        when "11110101110" => delta <= "000000111011111";
        when "11110101111" => delta <= "000000111011001";
        when "11110110000" => delta <= "000000111010100";
        when "11110110001" => delta <= "000000111001110";
        when "11110110010" => delta <= "000000111001000";
        when "11110110011" => delta <= "000000111000011";
        when "11110110100" => delta <= "000000110111101";
        when "11110110101" => delta <= "000000110110111";
        when "11110110110" => delta <= "000000110110010";
        when "11110110111" => delta <= "000000110101100";
        when "11110111000" => delta <= "000000110100111";
        when "11110111001" => delta <= "000000110100001";
        when "11110111010" => delta <= "000000110011011";
        when "11110111011" => delta <= "000000110010110";
        when "11110111100" => delta <= "000000110010000";
        when "11110111101" => delta <= "000000110001010";
        when "11110111110" => delta <= "000000110000101";
        when "11110111111" => delta <= "000000101111111";
        when "11111000000" => delta <= "000000101111001";
        when "11111000001" => delta <= "000000101110011";
        when "11111000010" => delta <= "000000101101110";
        when "11111000011" => delta <= "000000101101000";
        when "11111000100" => delta <= "000000101100010";
        when "11111000101" => delta <= "000000101011100";
        when "11111000110" => delta <= "000000101010111";
        when "11111000111" => delta <= "000000101010001";
        when "11111001000" => delta <= "000000101001011";
        when "11111001001" => delta <= "000000101000101";
        when "11111001010" => delta <= "000000101000000";
        when "11111001011" => delta <= "000000100111010";
        when "11111001100" => delta <= "000000100110100";
        when "11111001101" => delta <= "000000100101110";
        when "11111001110" => delta <= "000000100101000";
        when "11111001111" => delta <= "000000100100011";
        when "11111010000" => delta <= "000000100011101";
        when "11111010001" => delta <= "000000100010111";
        when "11111010010" => delta <= "000000100010001";
        when "11111010011" => delta <= "000000100001011";
        when "11111010100" => delta <= "000000100000101";
        when "11111010101" => delta <= "000000100000000";
        when "11111010110" => delta <= "000000011111010";
        when "11111010111" => delta <= "000000011110100";
        when "11111011000" => delta <= "000000011101110";
        when "11111011001" => delta <= "000000011101000";
        when "11111011010" => delta <= "000000011100010";
        when "11111011011" => delta <= "000000011011100";
        when "11111011100" => delta <= "000000011010110";
        when "11111011101" => delta <= "000000011010000";
        when "11111011110" => delta <= "000000011001011";
        when "11111011111" => delta <= "000000011000101";
        when "11111100000" => delta <= "000000010111111";
        when "11111100001" => delta <= "000000010111001";
        when "11111100010" => delta <= "000000010110011";
        when "11111100011" => delta <= "000000010101101";
        when "11111100100" => delta <= "000000010100111";
        when "11111100101" => delta <= "000000010100001";
        when "11111100110" => delta <= "000000010011011";
        when "11111100111" => delta <= "000000010010101";
        when "11111101000" => delta <= "000000010001111";
        when "11111101001" => delta <= "000000010001001";
        when "11111101010" => delta <= "000000010000011";
        when "11111101011" => delta <= "000000001111101";
        when "11111101100" => delta <= "000000001110111";
        when "11111101101" => delta <= "000000001110001";
        when "11111101110" => delta <= "000000001101011";
        when "11111101111" => delta <= "000000001100101";
        when "11111110000" => delta <= "000000001011111";
        when "11111110001" => delta <= "000000001011001";
        when "11111110010" => delta <= "000000001010010";
        when "11111110011" => delta <= "000000001001100";
        when "11111110100" => delta <= "000000001000110";
        when "11111110101" => delta <= "000000001000000";
        when "11111110110" => delta <= "000000000111010";
        when "11111110111" => delta <= "000000000110100";
        when "11111111000" => delta <= "000000000101110";
        when "11111111001" => delta <= "000000000101000";
        when "11111111010" => delta <= "000000000100010";
        when "11111111011" => delta <= "000000000011011";
        when "11111111100" => delta <= "000000000010101";
        when "11111111101" => delta <= "000000000001111";
        when "11111111110" => delta <= "000000000001001";
        when "11111111111" => delta <= "000000000000011";
    end case;
end process;

end Behavioral;
