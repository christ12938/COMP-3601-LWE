----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date: 11/16/2021 04:58:20 PM
-- Design Name:
-- Module Name: log_deltas - Behavioral
-- Project Name:
-- Target Devices:
-- Tool Versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE WORK.DATA_TYPES.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity exp_deltas is
    Port (frac : in unsigned(mE - 1 downto 0);
          delta : out unsigned(k_trunc-1 downto 0));
end exp_deltas;

architecture Behavioral of exp_deltas is
begin

process (frac)
begin
    case frac is
        when "000000000" => delta <= "000000000001001";
        when "000000001" => delta <= "000000000011101";
        when "000000010" => delta <= "000000000110000";
        when "000000011" => delta <= "000000001000100";
        when "000000100" => delta <= "000000001010111";
        when "000000101" => delta <= "000000001101010";
        when "000000110" => delta <= "000000001111110";
        when "000000111" => delta <= "000000010010001";
        when "000001000" => delta <= "000000010100100";
        when "000001001" => delta <= "000000010110111";
        when "000001010" => delta <= "000000011001010";
        when "000001011" => delta <= "000000011011101";
        when "000001100" => delta <= "000000011110000";
        when "000001101" => delta <= "000000100000011";
        when "000001110" => delta <= "000000100010110";
        when "000001111" => delta <= "000000100101000";
        when "000010000" => delta <= "000000100111011";
        when "000010001" => delta <= "000000101001110";
        when "000010010" => delta <= "000000101100000";
        when "000010011" => delta <= "000000101110011";
        when "000010100" => delta <= "000000110000101";
        when "000010101" => delta <= "000000110011000";
        when "000010110" => delta <= "000000110101010";
        when "000010111" => delta <= "000000110111100";
        when "000011000" => delta <= "000000111001110";
        when "000011001" => delta <= "000000111100000";
        when "000011010" => delta <= "000000111110010";
        when "000011011" => delta <= "000001000000100";
        when "000011100" => delta <= "000001000010110";
        when "000011101" => delta <= "000001000101000";
        when "000011110" => delta <= "000001000111010";
        when "000011111" => delta <= "000001001001100";
        when "000100000" => delta <= "000001001011101";
        when "000100001" => delta <= "000001001101111";
        when "000100010" => delta <= "000001010000001";
        when "000100011" => delta <= "000001010010010";
        when "000100100" => delta <= "000001010100011";
        when "000100101" => delta <= "000001010110101";
        when "000100110" => delta <= "000001011000110";
        when "000100111" => delta <= "000001011010111";
        when "000101000" => delta <= "000001011101001";
        when "000101001" => delta <= "000001011111010";
        when "000101010" => delta <= "000001100001011";
        when "000101011" => delta <= "000001100011100";
        when "000101100" => delta <= "000001100101101";
        when "000101101" => delta <= "000001100111101";
        when "000101110" => delta <= "000001101001110";
        when "000101111" => delta <= "000001101011111";
        when "000110000" => delta <= "000001101110000";
        when "000110001" => delta <= "000001110000000";
        when "000110010" => delta <= "000001110010001";
        when "000110011" => delta <= "000001110100001";
        when "000110100" => delta <= "000001110110010";
        when "000110101" => delta <= "000001111000010";
        when "000110110" => delta <= "000001111010010";
        when "000110111" => delta <= "000001111100010";
        when "000111000" => delta <= "000001111110011";
        when "000111001" => delta <= "000010000000011";
        when "000111010" => delta <= "000010000010011";
        when "000111011" => delta <= "000010000100011";
        when "000111100" => delta <= "000010000110011";
        when "000111101" => delta <= "000010001000010";
        when "000111110" => delta <= "000010001010010";
        when "000111111" => delta <= "000010001100010";
        when "001000000" => delta <= "000010001110001";
        when "001000001" => delta <= "000010010000001";
        when "001000010" => delta <= "000010010010000";
        when "001000011" => delta <= "000010010100000";
        when "001000100" => delta <= "000010010101111";
        when "001000101" => delta <= "000010010111111";
        when "001000110" => delta <= "000010011001110";
        when "001000111" => delta <= "000010011011101";
        when "001001000" => delta <= "000010011101100";
        when "001001001" => delta <= "000010011111011";
        when "001001010" => delta <= "000010100001010";
        when "001001011" => delta <= "000010100011001";
        when "001001100" => delta <= "000010100101000";
        when "001001101" => delta <= "000010100110111";
        when "001001110" => delta <= "000010101000101";
        when "001001111" => delta <= "000010101010100";
        when "001010000" => delta <= "000010101100010";
        when "001010001" => delta <= "000010101110001";
        when "001010010" => delta <= "000010101111111";
        when "001010011" => delta <= "000010110001110";
        when "001010100" => delta <= "000010110011100";
        when "001010101" => delta <= "000010110101010";
        when "001010110" => delta <= "000010110111000";
        when "001010111" => delta <= "000010111000111";
        when "001011000" => delta <= "000010111010101";
        when "001011001" => delta <= "000010111100010";
        when "001011010" => delta <= "000010111110000";
        when "001011011" => delta <= "000010111111110";
        when "001011100" => delta <= "000011000001100";
        when "001011101" => delta <= "000011000011010";
        when "001011110" => delta <= "000011000100111";
        when "001011111" => delta <= "000011000110101";
        when "001100000" => delta <= "000011001000010";
        when "001100001" => delta <= "000011001010000";
        when "001100010" => delta <= "000011001011101";
        when "001100011" => delta <= "000011001101010";
        when "001100100" => delta <= "000011001111000";
        when "001100101" => delta <= "000011010000101";
        when "001100110" => delta <= "000011010010010";
        when "001100111" => delta <= "000011010011111";
        when "001101000" => delta <= "000011010101100";
        when "001101001" => delta <= "000011010111001";
        when "001101010" => delta <= "000011011000101";
        when "001101011" => delta <= "000011011010010";
        when "001101100" => delta <= "000011011011111";
        when "001101101" => delta <= "000011011101011";
        when "001101110" => delta <= "000011011111000";
        when "001101111" => delta <= "000011100000100";
        when "001110000" => delta <= "000011100010001";
        when "001110001" => delta <= "000011100011101";
        when "001110010" => delta <= "000011100101001";
        when "001110011" => delta <= "000011100110101";
        when "001110100" => delta <= "000011101000001";
        when "001110101" => delta <= "000011101001101";
        when "001110110" => delta <= "000011101011001";
        when "001110111" => delta <= "000011101100101";
        when "001111000" => delta <= "000011101110001";
        when "001111001" => delta <= "000011101111101";
        when "001111010" => delta <= "000011110001001";
        when "001111011" => delta <= "000011110010100";
        when "001111100" => delta <= "000011110100000";
        when "001111101" => delta <= "000011110101011";
        when "001111110" => delta <= "000011110110111";
        when "001111111" => delta <= "000011111000010";
        when "010000000" => delta <= "000011111001101";
        when "010000001" => delta <= "000011111011000";
        when "010000010" => delta <= "000011111100011";
        when "010000011" => delta <= "000011111101110";
        when "010000100" => delta <= "000011111111001";
        when "010000101" => delta <= "000100000000100";
        when "010000110" => delta <= "000100000001111";
        when "010000111" => delta <= "000100000011010";
        when "010001000" => delta <= "000100000100100";
        when "010001001" => delta <= "000100000101111";
        when "010001010" => delta <= "000100000111010";
        when "010001011" => delta <= "000100001000100";
        when "010001100" => delta <= "000100001001110";
        when "010001101" => delta <= "000100001011001";
        when "010001110" => delta <= "000100001100011";
        when "010001111" => delta <= "000100001101101";
        when "010010000" => delta <= "000100001110111";
        when "010010001" => delta <= "000100010000001";
        when "010010010" => delta <= "000100010001011";
        when "010010011" => delta <= "000100010010101";
        when "010010100" => delta <= "000100010011111";
        when "010010101" => delta <= "000100010101001";
        when "010010110" => delta <= "000100010110010";
        when "010010111" => delta <= "000100010111100";
        when "010011000" => delta <= "000100011000101";
        when "010011001" => delta <= "000100011001111";
        when "010011010" => delta <= "000100011011000";
        when "010011011" => delta <= "000100011100001";
        when "010011100" => delta <= "000100011101011";
        when "010011101" => delta <= "000100011110100";
        when "010011110" => delta <= "000100011111101";
        when "010011111" => delta <= "000100100000110";
        when "010100000" => delta <= "000100100001111";
        when "010100001" => delta <= "000100100011000";
        when "010100010" => delta <= "000100100100000";
        when "010100011" => delta <= "000100100101001";
        when "010100100" => delta <= "000100100110010";
        when "010100101" => delta <= "000100100111010";
        when "010100110" => delta <= "000100101000011";
        when "010100111" => delta <= "000100101001011";
        when "010101000" => delta <= "000100101010011";
        when "010101001" => delta <= "000100101011011";
        when "010101010" => delta <= "000100101100100";
        when "010101011" => delta <= "000100101101100";
        when "010101100" => delta <= "000100101110100";
        when "010101101" => delta <= "000100101111100";
        when "010101110" => delta <= "000100110000100";
        when "010101111" => delta <= "000100110001011";
        when "010110000" => delta <= "000100110010011";
        when "010110001" => delta <= "000100110011011";
        when "010110010" => delta <= "000100110100010";
        when "010110011" => delta <= "000100110101010";
        when "010110100" => delta <= "000100110110001";
        when "010110101" => delta <= "000100110111000";
        when "010110110" => delta <= "000100111000000";
        when "010110111" => delta <= "000100111000111";
        when "010111000" => delta <= "000100111001110";
        when "010111001" => delta <= "000100111010101";
        when "010111010" => delta <= "000100111011100";
        when "010111011" => delta <= "000100111100011";
        when "010111100" => delta <= "000100111101001";
        when "010111101" => delta <= "000100111110000";
        when "010111110" => delta <= "000100111110111";
        when "010111111" => delta <= "000100111111101";
        when "011000000" => delta <= "000101000000100";
        when "011000001" => delta <= "000101000001010";
        when "011000010" => delta <= "000101000010001";
        when "011000011" => delta <= "000101000010111";
        when "011000100" => delta <= "000101000011101";
        when "011000101" => delta <= "000101000100011";
        when "011000110" => delta <= "000101000101001";
        when "011000111" => delta <= "000101000101111";
        when "011001000" => delta <= "000101000110101";
        when "011001001" => delta <= "000101000111011";
        when "011001010" => delta <= "000101001000000";
        when "011001011" => delta <= "000101001000110";
        when "011001100" => delta <= "000101001001011";
        when "011001101" => delta <= "000101001010001";
        when "011001110" => delta <= "000101001010110";
        when "011001111" => delta <= "000101001011011";
        when "011010000" => delta <= "000101001100001";
        when "011010001" => delta <= "000101001100110";
        when "011010010" => delta <= "000101001101011";
        when "011010011" => delta <= "000101001110000";
        when "011010100" => delta <= "000101001110101";
        when "011010101" => delta <= "000101001111010";
        when "011010110" => delta <= "000101001111110";
        when "011010111" => delta <= "000101010000011";
        when "011011000" => delta <= "000101010001000";
        when "011011001" => delta <= "000101010001100";
        when "011011010" => delta <= "000101010010000";
        when "011011011" => delta <= "000101010010101";
        when "011011100" => delta <= "000101010011001";
        when "011011101" => delta <= "000101010011101";
        when "011011110" => delta <= "000101010100001";
        when "011011111" => delta <= "000101010100101";
        when "011100000" => delta <= "000101010101001";
        when "011100001" => delta <= "000101010101101";
        when "011100010" => delta <= "000101010110001";
        when "011100011" => delta <= "000101010110100";
        when "011100100" => delta <= "000101010111000";
        when "011100101" => delta <= "000101010111100";
        when "011100110" => delta <= "000101010111111";
        when "011100111" => delta <= "000101011000010";
        when "011101000" => delta <= "000101011000110";
        when "011101001" => delta <= "000101011001001";
        when "011101010" => delta <= "000101011001100";
        when "011101011" => delta <= "000101011001111";
        when "011101100" => delta <= "000101011010010";
        when "011101101" => delta <= "000101011010101";
        when "011101110" => delta <= "000101011011000";
        when "011101111" => delta <= "000101011011010";
        when "011110000" => delta <= "000101011011101";
        when "011110001" => delta <= "000101011011111";
        when "011110010" => delta <= "000101011100010";
        when "011110011" => delta <= "000101011100100";
        when "011110100" => delta <= "000101011100110";
        when "011110101" => delta <= "000101011101001";
        when "011110110" => delta <= "000101011101011";
        when "011110111" => delta <= "000101011101101";
        when "011111000" => delta <= "000101011101111";
        when "011111001" => delta <= "000101011110001";
        when "011111010" => delta <= "000101011110010";
        when "011111011" => delta <= "000101011110100";
        when "011111100" => delta <= "000101011110110";
        when "011111101" => delta <= "000101011110111";
        when "011111110" => delta <= "000101011111001";
        when "011111111" => delta <= "000101011111010";
        when "100000000" => delta <= "000101011111011";
        when "100000001" => delta <= "000101011111100";
        when "100000010" => delta <= "000101011111101";
        when "100000011" => delta <= "000101011111110";
        when "100000100" => delta <= "000101011111111";
        when "100000101" => delta <= "000101100000000";
        when "100000110" => delta <= "000101100000001";
        when "100000111" => delta <= "000101100000010";
        when "100001000" => delta <= "000101100000010";
        when "100001001" => delta <= "000101100000011";
        when "100001010" => delta <= "000101100000011";
        when "100001011" => delta <= "000101100000011";
        when "100001100" => delta <= "000101100000100";
        when "100001101" => delta <= "000101100000100";
        when "100001110" => delta <= "000101100000100";
        when "100001111" => delta <= "000101100000100";
        when "100010000" => delta <= "000101100000100";
        when "100010001" => delta <= "000101100000100";
        when "100010010" => delta <= "000101100000011";
        when "100010011" => delta <= "000101100000011";
        when "100010100" => delta <= "000101100000010";
        when "100010101" => delta <= "000101100000010";
        when "100010110" => delta <= "000101100000001";
        when "100010111" => delta <= "000101100000001";
        when "100011000" => delta <= "000101100000000";
        when "100011001" => delta <= "000101011111111";
        when "100011010" => delta <= "000101011111110";
        when "100011011" => delta <= "000101011111101";
        when "100011100" => delta <= "000101011111100";
        when "100011101" => delta <= "000101011111010";
        when "100011110" => delta <= "000101011111001";
        when "100011111" => delta <= "000101011111000";
        when "100100000" => delta <= "000101011110110";
        when "100100001" => delta <= "000101011110100";
        when "100100010" => delta <= "000101011110011";
        when "100100011" => delta <= "000101011110001";
        when "100100100" => delta <= "000101011101111";
        when "100100101" => delta <= "000101011101101";
        when "100100110" => delta <= "000101011101011";
        when "100100111" => delta <= "000101011101001";
        when "100101000" => delta <= "000101011100111";
        when "100101001" => delta <= "000101011100100";
        when "100101010" => delta <= "000101011100010";
        when "100101011" => delta <= "000101011100000";
        when "100101100" => delta <= "000101011011101";
        when "100101101" => delta <= "000101011011010";
        when "100101110" => delta <= "000101011011000";
        when "100101111" => delta <= "000101011010101";
        when "100110000" => delta <= "000101011010010";
        when "100110001" => delta <= "000101011001111";
        when "100110010" => delta <= "000101011001100";
        when "100110011" => delta <= "000101011001000";
        when "100110100" => delta <= "000101011000101";
        when "100110101" => delta <= "000101011000010";
        when "100110110" => delta <= "000101010111110";
        when "100110111" => delta <= "000101010111011";
        when "100111000" => delta <= "000101010110111";
        when "100111001" => delta <= "000101010110011";
        when "100111010" => delta <= "000101010101111";
        when "100111011" => delta <= "000101010101011";
        when "100111100" => delta <= "000101010100111";
        when "100111101" => delta <= "000101010100011";
        when "100111110" => delta <= "000101010011111";
        when "100111111" => delta <= "000101010011011";
        when "101000000" => delta <= "000101010010110";
        when "101000001" => delta <= "000101010010010";
        when "101000010" => delta <= "000101010001101";
        when "101000011" => delta <= "000101010001000";
        when "101000100" => delta <= "000101010000100";
        when "101000101" => delta <= "000101001111111";
        when "101000110" => delta <= "000101001111010";
        when "101000111" => delta <= "000101001110101";
        when "101001000" => delta <= "000101001101111";
        when "101001001" => delta <= "000101001101010";
        when "101001010" => delta <= "000101001100101";
        when "101001011" => delta <= "000101001011111";
        when "101001100" => delta <= "000101001011010";
        when "101001101" => delta <= "000101001010100";
        when "101001110" => delta <= "000101001001111";
        when "101001111" => delta <= "000101001001001";
        when "101010000" => delta <= "000101001000011";
        when "101010001" => delta <= "000101000111101";
        when "101010010" => delta <= "000101000110111";
        when "101010011" => delta <= "000101000110001";
        when "101010100" => delta <= "000101000101010";
        when "101010101" => delta <= "000101000100100";
        when "101010110" => delta <= "000101000011101";
        when "101010111" => delta <= "000101000010111";
        when "101011000" => delta <= "000101000010000";
        when "101011001" => delta <= "000101000001001";
        when "101011010" => delta <= "000101000000010";
        when "101011011" => delta <= "000100111111100";
        when "101011100" => delta <= "000100111110100";
        when "101011101" => delta <= "000100111101101";
        when "101011110" => delta <= "000100111100110";
        when "101011111" => delta <= "000100111011111";
        when "101100000" => delta <= "000100111010111";
        when "101100001" => delta <= "000100111010000";
        when "101100010" => delta <= "000100111001000";
        when "101100011" => delta <= "000100111000000";
        when "101100100" => delta <= "000100110111001";
        when "101100101" => delta <= "000100110110001";
        when "101100110" => delta <= "000100110101001";
        when "101100111" => delta <= "000100110100000";
        when "101101000" => delta <= "000100110011000";
        when "101101001" => delta <= "000100110010000";
        when "101101010" => delta <= "000100110000111";
        when "101101011" => delta <= "000100101111111";
        when "101101100" => delta <= "000100101110110";
        when "101101101" => delta <= "000100101101110";
        when "101101110" => delta <= "000100101100101";
        when "101101111" => delta <= "000100101011100";
        when "101110000" => delta <= "000100101010011";
        when "101110001" => delta <= "000100101001010";
        when "101110010" => delta <= "000100101000001";
        when "101110011" => delta <= "000100100110111";
        when "101110100" => delta <= "000100100101110";
        when "101110101" => delta <= "000100100100100";
        when "101110110" => delta <= "000100100011011";
        when "101110111" => delta <= "000100100010001";
        when "101111000" => delta <= "000100100000111";
        when "101111001" => delta <= "000100011111101";
        when "101111010" => delta <= "000100011110011";
        when "101111011" => delta <= "000100011101001";
        when "101111100" => delta <= "000100011011111";
        when "101111101" => delta <= "000100011010101";
        when "101111110" => delta <= "000100011001010";
        when "101111111" => delta <= "000100011000000";
        when "110000000" => delta <= "000100010110101";
        when "110000001" => delta <= "000100010101011";
        when "110000010" => delta <= "000100010100000";
        when "110000011" => delta <= "000100010010101";
        when "110000100" => delta <= "000100010001010";
        when "110000101" => delta <= "000100001111111";
        when "110000110" => delta <= "000100001110100";
        when "110000111" => delta <= "000100001101000";
        when "110001000" => delta <= "000100001011101";
        when "110001001" => delta <= "000100001010001";
        when "110001010" => delta <= "000100001000110";
        when "110001011" => delta <= "000100000111010";
        when "110001100" => delta <= "000100000101110";
        when "110001101" => delta <= "000100000100010";
        when "110001110" => delta <= "000100000010110";
        when "110001111" => delta <= "000100000001010";
        when "110010000" => delta <= "000011111111110";
        when "110010001" => delta <= "000011111110001";
        when "110010010" => delta <= "000011111100101";
        when "110010011" => delta <= "000011111011000";
        when "110010100" => delta <= "000011111001100";
        when "110010101" => delta <= "000011110111111";
        when "110010110" => delta <= "000011110110010";
        when "110010111" => delta <= "000011110100101";
        when "110011000" => delta <= "000011110011000";
        when "110011001" => delta <= "000011110001011";
        when "110011010" => delta <= "000011101111110";
        when "110011011" => delta <= "000011101110000";
        when "110011100" => delta <= "000011101100011";
        when "110011101" => delta <= "000011101010101";
        when "110011110" => delta <= "000011101000111";
        when "110011111" => delta <= "000011100111010";
        when "110100000" => delta <= "000011100101100";
        when "110100001" => delta <= "000011100011110";
        when "110100010" => delta <= "000011100010000";
        when "110100011" => delta <= "000011100000001";
        when "110100100" => delta <= "000011011110011";
        when "110100101" => delta <= "000011011100101";
        when "110100110" => delta <= "000011011010110";
        when "110100111" => delta <= "000011011000111";
        when "110101000" => delta <= "000011010111001";
        when "110101001" => delta <= "000011010101010";
        when "110101010" => delta <= "000011010011011";
        when "110101011" => delta <= "000011010001100";
        when "110101100" => delta <= "000011001111101";
        when "110101101" => delta <= "000011001101101";
        when "110101110" => delta <= "000011001011110";
        when "110101111" => delta <= "000011001001110";
        when "110110000" => delta <= "000011000111111";
        when "110110001" => delta <= "000011000101111";
        when "110110010" => delta <= "000011000011111";
        when "110110011" => delta <= "000011000001111";
        when "110110100" => delta <= "000010111111111";
        when "110110101" => delta <= "000010111101111";
        when "110110110" => delta <= "000010111011111";
        when "110110111" => delta <= "000010111001110";
        when "110111000" => delta <= "000010110111110";
        when "110111001" => delta <= "000010110101101";
        when "110111010" => delta <= "000010110011101";
        when "110111011" => delta <= "000010110001100";
        when "110111100" => delta <= "000010101111011";
        when "110111101" => delta <= "000010101101010";
        when "110111110" => delta <= "000010101011001";
        when "110111111" => delta <= "000010101001000";
        when "111000000" => delta <= "000010100110110";
        when "111000001" => delta <= "000010100100101";
        when "111000010" => delta <= "000010100010011";
        when "111000011" => delta <= "000010100000001";
        when "111000100" => delta <= "000010011110000";
        when "111000101" => delta <= "000010011011110";
        when "111000110" => delta <= "000010011001100";
        when "111000111" => delta <= "000010010111010";
        when "111001000" => delta <= "000010010100111";
        when "111001001" => delta <= "000010010010101";
        when "111001010" => delta <= "000010010000010";
        when "111001011" => delta <= "000010001110000";
        when "111001100" => delta <= "000010001011101";
        when "111001101" => delta <= "000010001001010";
        when "111001110" => delta <= "000010000111000";
        when "111001111" => delta <= "000010000100100";
        when "111010000" => delta <= "000010000010001";
        when "111010001" => delta <= "000001111111110";
        when "111010010" => delta <= "000001111101011";
        when "111010011" => delta <= "000001111010111";
        when "111010100" => delta <= "000001111000100";
        when "111010101" => delta <= "000001110110000";
        when "111010110" => delta <= "000001110011100";
        when "111010111" => delta <= "000001110001000";
        when "111011000" => delta <= "000001101110100";
        when "111011001" => delta <= "000001101100000";
        when "111011010" => delta <= "000001101001100";
        when "111011011" => delta <= "000001100110111";
        when "111011100" => delta <= "000001100100011";
        when "111011101" => delta <= "000001100001110";
        when "111011110" => delta <= "000001011111001";
        when "111011111" => delta <= "000001011100101";
        when "111100000" => delta <= "000001011010000";
        when "111100001" => delta <= "000001010111011";
        when "111100010" => delta <= "000001010100101";
        when "111100011" => delta <= "000001010010000";
        when "111100100" => delta <= "000001001111011";
        when "111100101" => delta <= "000001001100101";
        when "111100110" => delta <= "000001001001111";
        when "111100111" => delta <= "000001000111010";
        when "111101000" => delta <= "000001000100100";
        when "111101001" => delta <= "000001000001110";
        when "111101010" => delta <= "000000111111000";
        when "111101011" => delta <= "000000111100001";
        when "111101100" => delta <= "000000111001011";
        when "111101101" => delta <= "000000110110101";
        when "111101110" => delta <= "000000110011110";
        when "111101111" => delta <= "000000110000111";
        when "111110000" => delta <= "000000101110001";
        when "111110001" => delta <= "000000101011010";
        when "111110010" => delta <= "000000101000011";
        when "111110011" => delta <= "000000100101011";
        when "111110100" => delta <= "000000100010100";
        when "111110101" => delta <= "000000011111101";
        when "111110110" => delta <= "000000011100101";
        when "111110111" => delta <= "000000011001110";
        when "111111000" => delta <= "000000010110110";
        when "111111001" => delta <= "000000010011110";
        when "111111010" => delta <= "000000010000110";
        when "111111011" => delta <= "000000001101110";
        when "111111100" => delta <= "000000001010101";
        when "111111101" => delta <= "000000000111101";
        when "111111110" => delta <= "000000000100101";
        when "111111111" => delta <= "000000000001100";
        when others => delta <= "000000000000000";

    end case;
end process;

end Behavioral;
